LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY rom IS
  PORT (
    address : IN STD_ULOGIC_VECTOR(14 DOWNTO 0);
    data_out : OUT STD_ULOGIC_VECTOR(15 DOWNTO 0));
END ENTITY;

ARCHITECTURE behavioural OF rom IS
  TYPE ROM_type IS ARRAY (0 TO 32767) OF STD_ULOGIC_VECTOR(15 DOWNTO 0);
  CONSTANT ROM : ROM_type := (0 => "1001101111100101", 1 => "0000011110011111", 2 => "1001111000000011", 3 => "0101000011010100", 4 => "1000011100011111", 5 => "1010011111011011", 6 => "0001011101010111", 7 => "1111101011100011", 8 => "1010110101000001", 9 => "1011111011011110", 10 => "0100000101111000", 11 => "1111111011000111", 12 => "1111001100010100", 13 => "0110101000001111", 14 => "1100010010000010", 15 => "1110000010101110", 16 => "0100011100101101", 17 => "0001111011110110", 18 => "1000110001010010", 19 => "0110011100100110", 20 => "0001010000011101", 21 => "0000001111111110", 22 => "1010101010111101", 23 => "1010010001011010", 24 => "1100001001101101", 25 => "1000111100100111", 26 => "0010010010111010", 27 => "0111001011001011", 28 => "1011000011101111", 29 => "0111101010000001", 30 => "1000100111110111", 31 => "1111100111001100", 32 => "0011101110000010", 33 => "1010001000101001", 34 => "0110010010010000", 35 => "1000100000010001", 36 => "0100101010101011", 37 => "1011010101001001", 38 => "0001101110001001", 39 => "0101001110101000", 40 => "1001010110010110", 41 => "1011000100000100", 42 => "0000001010101000", 43 => "1011011100101000", 44 => "1110100000111111", 45 => "0001110000010000", 46 => "0110000110101010", 47 => "1110010011100011", 48 => "0001000111110010", 49 => "1010011111100001", 50 => "0000010000011100", 51 => "1001110111110010", 52 => "0010010100010111", 53 => "0011110101110101", 54 => "1001110101000111", 55 => "1111100100101101", 56 => "1000010110001100", 57 => "0010111000010001", 58 => "0011111011011101", 59 => "1110000101101010", 60 => "1111101000011100", 61 => "1010110000100001", 62 => "1100111001001111", 63 => "1000010010010100", 64 => "1111111011100000", 65 => "0011011110000101", 66 => "1111011111011101", 67 => "0101101100101011", 68 => "0110010100100010", 69 => "0101101000001111", 70 => "1100101001010111", 71 => "0011010101100100", 72 => "0101110001110001", 73 => "0100000111010001", 74 => "1011011011010011", 75 => "0011000000000111", 76 => "1001100111010111", 77 => "0100001101110110", 78 => "1101001010011110", 79 => "0011000001110100", 80 => "1011111100010010", 81 => "1001000001111111", 82 => "0000001100111001", 83 => "1011010011111111", 84 => "0100010110111001", 85 => "0101110001000001", 86 => "1100111011000000", 87 => "1101010000001110", 88 => "0100111101011100", 89 => "1000111010010111", 90 => "0000111110011110", 91 => "1011001001111101", 92 => "1110100010100110", 93 => "0110010111110110", 94 => "0111111101000011", 95 => "0110001110110101", 96 => "0111110110101001", 97 => "0011000110001000", 98 => "0100001011011001", 99 => "0011100010100001", 100 => "1111110100110111", 101 => "1101010101100111", 102 => "0001001101101110", 103 => "0110101111101000", 104 => "1010001110011111", 105 => "1011100000011001", 106 => "0011100011111000", 107 => "1101011001100011", 108 => "0110101110101001", 109 => "0110011001011010", 110 => "0101100011100101", 111 => "0111001100010001", 112 => "1101101011110111", 113 => "0110111101100010", 114 => "0000110101001001", 115 => "1100110100100000", 116 => "0011101011010000", 117 => "0110110110010001", 118 => "0001110010011101", 119 => "1000011010101011", 120 => "0100011100001000", 121 => "0100011000001100", 122 => "1000001100001000", 123 => "1010000100100101", 124 => "0100101101100000", 125 => "1011110100110010", 126 => "0111101100101101", 127 => "1100001000011010", 128 => "0100110000011001", 129 => "1000011110010000", 130 => "1100110110111000", 131 => "0101110010010011", 132 => "0000110100000010", 133 => "1010101100001000", 134 => "1101111101010010", 135 => "0001001010010011", 136 => "0001110101010110", 137 => "1010111101111011", 138 => "0000010000101000", 139 => "1010001110111101", 140 => "1010100011101100", 141 => "0011100010000111", 142 => "1000001011110100", 143 => "0101001100000011", 144 => "1010011111010011", 145 => "1111011000001001", 146 => "0011011111010011", 147 => "1101111100010100", 148 => "0101101011001111", 149 => "0011000110001110", 150 => "1101111010010101", 151 => "1101100110000011", 152 => "1000000110110110", 153 => "0000010000100111", 154 => "0101010100011111", 155 => "0001010001100101", 156 => "1011101011100011", 157 => "1000110000010101", 158 => "1101001110101001", 159 => "0101100101011011", 160 => "0001111001100100", 161 => "1101011110011001", 162 => "1001011111100101", 163 => "1000010010110101", 164 => "0001100010000011", 165 => "1110111001111111", 166 => "1100111010101100", 167 => "0011011100011110", 168 => "0110001111100101", 169 => "1000000101100000", 170 => "1101101001000111", 171 => "1100101011111010", 172 => "1110001010110000", 173 => "1011000010011111", 174 => "1001100110101111", 175 => "0111011110011001", 176 => "0110000000101001", 177 => "1101001101000010", 178 => "1011101111001001", 179 => "0101110110101101", 180 => "1011001101011011", 181 => "1100110010110011", 182 => "1001011001000000", 183 => "0101001001101100", 184 => "1100101101110001", 185 => "1000000100001111", 186 => "0001110011101110", 187 => "0001001111001111", 188 => "0100011110001000", 189 => "0100011100111010", 190 => "1100000010010111", 191 => "1101110011001100", 192 => "1011100111011100", 193 => "1010011011101000", 194 => "0000010110100111", 195 => "0100111100011010", 196 => "0110011001000001", 197 => "0010010011100010", 198 => "0100000100010011", 199 => "0011111111000010", 200 => "1000010110101010", 201 => "0011111101010001", 202 => "1000100010010110", 203 => "0111011100000100", 204 => "1101000010101011", 205 => "1111001000100110", 206 => "0001101100010011", 207 => "1000110110101001", 208 => "0000010110000101", 209 => "0110100011100000", 210 => "1001011000000000", 211 => "1111110111100101", 212 => "0010011010101111", 213 => "1001111011000010", 214 => "1001010101011011", 215 => "0110001111110000", 216 => "0001111111010000", 217 => "1110001100101010", 218 => "0011001011001011", 219 => "0100110001000100", 220 => "1010000010110011", 221 => "1010111111111011", 222 => "1101011000010001", 223 => "1010100001111010", 224 => "0101011001101010", 225 => "1111100111001100", 226 => "1010010111101110", 227 => "1100110010011110", 228 => "1001110011000101", 229 => "0000101100110010", 230 => "1111000001110110", 231 => "1001011001110110", 232 => "0110110011010101", 233 => "0000011011000101", 234 => "0011011001000100", 235 => "0111000111110010", 236 => "0110100101100010", 237 => "1101011010100111", 238 => "0001100111100110", 239 => "0101100111101100", 240 => "1011111010101101", 241 => "0101101011110100", 242 => "0100011001110110", 243 => "1010010110010100", 244 => "0001100011101001", 245 => "1011110000000001", 246 => "0001110000010101", 247 => "1101010110100101", 248 => "1111111011101101", 249 => "1100011000100110", 250 => "1100011011000101", 251 => "1101000010011011", 252 => "0110001011011110", 253 => "0011010010001110", 254 => "1100100100001110", 255 => "0000110000111001", 256 => "0011111111101110", 257 => "1100011000010011", 258 => "0100010110110100", 259 => "1001111111101000", 260 => "0101000110111110", 261 => "1100111100100100", 262 => "1011000000011100", 263 => "0111100010001000", 264 => "1111110111101111", 265 => "1111100100010011", 266 => "1100001011001101", 267 => "0001111001101100", 268 => "0111001000010001", 269 => "0100111010001010", 270 => "0011111110111100", 271 => "1011100100000000", 272 => "1001100110011101", 273 => "0000010110110001", 274 => "1101100011011110", 275 => "1111101011110111", 276 => "0010001111100100", 277 => "1001111011100011", 278 => "1000101111101000", 279 => "1100000100110000", 280 => "1110001111010000", 281 => "0100011010000111", 282 => "1010111111001010", 283 => "0111010010010000", 284 => "0000011000111100", 285 => "1010111001000011", 286 => "1010101000000100", 287 => "0010001000100010", 288 => "1111101100110011", 289 => "1100000101000000", 290 => "0000011110011101", 291 => "1000010011101000", 292 => "1100000111001110", 293 => "1000011000001010", 294 => "1000001111110101", 295 => "1011010000101000", 296 => "1100101110101100", 297 => "1010101100100010", 298 => "0001011010110110", 299 => "0001011010000111", 300 => "0110111111011101", 301 => "0101111001010001", 302 => "0100000001111011", 303 => "0001001110101111", 304 => "1101000001010001", 305 => "1011100010100001", 306 => "1001101011111101", 307 => "1100011011010100", 308 => "0001001100000101", 309 => "1110000010110100", 310 => "0100101110001101", 311 => "0010001010010011", 312 => "1101001001000010", 313 => "1101011110111010", 314 => "1100000011000100", 315 => "1011010001001100", 316 => "0011100000000011", 317 => "1100110000000101", 318 => "1011001001110101", 319 => "1111011001100010", 320 => "1101100000001110", 321 => "0001001101011100", 322 => "1010101011101110", 323 => "0100000000101001", 324 => "1101010000100110", 325 => "1010111011111110", 326 => "1011101100010000", 327 => "1011011111110000", 328 => "1011100110011011", 329 => "1101001111001001", 330 => "1111110010101000", 331 => "1111100010010001", 332 => "0111100100000111", 333 => "0010111100000111", 334 => "0111000100010111", 335 => "0011111001111001", 336 => "1100010010010100", 337 => "0001101001000010", 338 => "0011010100101010", 339 => "1000110100101011", 340 => "0100100111010111", 341 => "0101101101001110", 342 => "0011111011000110", 343 => "1101100101000010", 344 => "1011000010001111", 345 => "0010001101111101", 346 => "1111010101101011", 347 => "1111101100100010", 348 => "0101101000001100", 349 => "0100010100111010", 350 => "1001100110110010", 351 => "0101111111001110", 352 => "1100001001000111", 353 => "1001001101101001", 354 => "1001101010110000", 355 => "1010100111111101", 356 => "1011011110101011", 357 => "0010001110101110", 358 => "1100000110101010", 359 => "1001110010101000", 360 => "1111010100101011", 361 => "0001011001001000", 362 => "0011101000111111", 363 => "0110110010011100", 364 => "0011110010100010", 365 => "1000010100110100", 366 => "1000010000011100", 367 => "1101011111110110", 368 => "1000011100110100", 369 => "1101100110110010", 370 => "0110011100110011", 371 => "0011011111011100", 372 => "1111011011100000", 373 => "0111000000011111", 374 => "0000110001101010", 375 => "1011000111100010", 376 => "0010001011100001", 377 => "1011010110111101", 378 => "0000111101100111", 379 => "1110101111000011", 380 => "1000010011111011", 381 => "0001111100111011", 382 => "0100001101110010", 383 => "0100001110101001", 384 => "0001010010111001", 385 => "0010011101000101", 386 => "1011100111101110", 387 => "1000011011110110", 388 => "1011101101111111", 389 => "0100011011000111", 390 => "1111110110010111", 391 => "1111111000101010", 392 => "0001011001100100", 393 => "1100111111000011", 394 => "0000110001000110", 395 => "0010001010100011", 396 => "1100001000110100", 397 => "1001100001000101", 398 => "0001001101111101", 399 => "0101101001101100", 400 => "0000100010010001", 401 => "0011011000001011", 402 => "1011111110111101", 403 => "1100001100011011", 404 => "0110011111110010", 405 => "0111100110100010", 406 => "0110110100101000", 407 => "1100100100001101", 408 => "0001110110110111", 409 => "1001010000111010", 410 => "1010000101100000", 411 => "0111100111111000", 412 => "1110110100100000", 413 => "0000111011110011", 414 => "1111100000101111", 415 => "1010000100001010", 416 => "1101101011000010", 417 => "1001011101100100", 418 => "1000010100011001", 419 => "0110000000101101", 420 => "1111001100100000", 421 => "1101010101000011", 422 => "1001010010000111", 423 => "1110110101100000", 424 => "1101100010100111", 425 => "0110101101000000", 426 => "1101111010000110", 427 => "1100000110001001", 428 => "1000101100011110", 429 => "1110100110100101", 430 => "1101110011000000", 431 => "1010111110010110", 432 => "0101101100111001", 433 => "1011010100001010", 434 => "1011001001110000", 435 => "1001110101011101", 436 => "0011011001010110", 437 => "0011100111001111", 438 => "1000101100001001", 439 => "0000010000011001", 440 => "0101001100101010", 441 => "1101001111010101", 442 => "1100110010100110", 443 => "0001100001011100", 444 => "0000010010110110", 445 => "1001010111011111", 446 => "1011101010001110", 447 => "1011001000100101", 448 => "1000111000001011", 449 => "0000001101000111", 450 => "0111001000010001", 451 => "0001110111010111", 452 => "0000101011001000", 453 => "1011000000010010", 454 => "1111111011101001", 455 => "1011011001111001", 456 => "0010001110011001", 457 => "0001011111010110", 458 => "0101000100111111", 459 => "1001010111100100", 460 => "1110011000101000", 461 => "1010110011110011", 462 => "0100101011011111", 463 => "0000110011110100", 464 => "0100100101111011", 465 => "0001100101101011", 466 => "0101011011001100", 467 => "0100110101111110", 468 => "1010111101101011", 469 => "0011001100100000", 470 => "1001110001111100", 471 => "1101100111010110", 472 => "1000011111111010", 473 => "1011000011110000", 474 => "1001000100110110", 475 => "0101000001111110", 476 => "1110110111110011", 477 => "1101000100010011", 478 => "1110010101010110", 479 => "0001111111011110", 480 => "0110110000100010", 481 => "1001110001100111", 482 => "1010000111010100", 483 => "0010110100110110", 484 => "1111000001101100", 485 => "0010110000101001", 486 => "1000010000110010", 487 => "0001111010111010", 488 => "1011100000101100", 489 => "1111000101101110", 490 => "0100010111011001", 491 => "1010111110010111", 492 => "1101000011000101", 493 => "0000111110011010", 494 => "0111110011111000", 495 => "0010010001010101", 496 => "1011100000001111", 497 => "1100000111100100", 498 => "1001011010110101", 499 => "0000111000011101", 500 => "0001101001010101", 501 => "0000011110110001", 502 => "1101110110101100", 503 => "0110101111100000", 504 => "1001000000110011", 505 => "1011011001001101", 506 => "1001000100101101", 507 => "0100000010011011", 508 => "0000000111111011", 509 => "0101111111000001", 510 => "0111110010010000", 511 => "1101010110100011", 512 => "0000100111100110", 513 => "0001100101010000", 514 => "0000011000001111", 515 => "0100010100001101", 516 => "1010111001100001", 517 => "0001001110111100", 518 => "1110001000101100", 519 => "1110010011001010", 520 => "0110010111100010", 521 => "1111001101100011", 522 => "0010000011001101", 523 => "0001000111100100", 524 => "0001110100100000", 525 => "1111110111110100", 526 => "0000110010111100", 527 => "0111000111000000", 528 => "0110111010011111", 529 => "1111000101111010", 530 => "0011101001110010", 531 => "0101000001100000", 532 => "1110000011011100", 533 => "1001101101100100", 534 => "0101111110100111", 535 => "1101111001100100", 536 => "1111100011100011", 537 => "0110111111101111", 538 => "1101011011101011", 539 => "1110110000100000", 540 => "0101000100010001", 541 => "0001010100110111", 542 => "1000000101110110", 543 => "0100111111011001", 544 => "1110110010100100", 545 => "0110101100101011", 546 => "1001010101011011", 547 => "1010110000100101", 548 => "1000101111000101", 549 => "0001111100101000", 550 => "1010011001001110", 551 => "1100100000111101", 552 => "1101000011010001", 553 => "1111101001101100", 554 => "1110100010011100", 555 => "0001101110011111", 556 => "1000000001111100", 557 => "1111110001110000", 558 => "1000110011010001", 559 => "1101101111111111", 560 => "0111110111100110", 561 => "0111101001000111", 562 => "0011111101000011", 563 => "1101001100110101", 564 => "1111011110011111", 565 => "0000001100100001", 566 => "1111111110111000", 567 => "0010101000101100", 568 => "0110010110010101", 569 => "1111110110101111", 570 => "0010011100000011", 571 => "1110011100100010", 572 => "0000111011111010", 573 => "1000111010100000", 574 => "1000000110010010", 575 => "0101100010010111", 576 => "1000000011101001", 577 => "0010110011110011", 578 => "1101011111000100", 579 => "0101000011110100", 580 => "1100111100000110", 581 => "1001011101011111", 582 => "0010011111010011", 583 => "1100000101010010", 584 => "1010101111010000", 585 => "1110000000001001", 586 => "0011111011111101", 587 => "0100011100011110", 588 => "1010101100101010", 589 => "0111111001010101", 590 => "1010101011000011", 591 => "0110110011100101", 592 => "0100001110110001", 593 => "1000110011100110", 594 => "0000000110010100", 595 => "0010110100011011", 596 => "0010011111000111", 597 => "1101010110100111", 598 => "1101100100101001", 599 => "0011001100110010", 600 => "1100011110011000", 601 => "0101111111010111", 602 => "1100110001110000", 603 => "1100010111110101", 604 => "1111111001101101", 605 => "1101101100011001", 606 => "1011001110101110", 607 => "0010001100111101", 608 => "1100111011110101", 609 => "0000010111010101", 610 => "1011000111101011", 611 => "1111101001110111", 612 => "0011101001011100", 613 => "0000000011111010", 614 => "0000010110110100", 615 => "0001000111110100", 616 => "1011010010011010", 617 => "1101100001001000", 618 => "0111010001100110", 619 => "1111001110010011", 620 => "0110011111001000", 621 => "0000001010111110", 622 => "1101111010000000", 623 => "1110001101101001", 624 => "0010101111001000", 625 => "1111111010010010", 626 => "0001000111000011", 627 => "1110110100001011", 628 => "1011000001101001", 629 => "1101101100110011", 630 => "0110100100100011", 631 => "0111100100011001", 632 => "1110110101111101", 633 => "1111110101101110", 634 => "1010111000010100", 635 => "1000001010111010", 636 => "0101100011101100", 637 => "1110000010000010", 638 => "0010000001001000", 639 => "0111110000010011", 640 => "1000010000100111", 641 => "1101110001000100", 642 => "0101010000110010", 643 => "0001010001000010", 644 => "0000111100000000", 645 => "1010011001010110", 646 => "1010101001101100", 647 => "1101110100011000", 648 => "0101000010011110", 649 => "1111010001100100", 650 => "1000000101001011", 651 => "1001011101111100", 652 => "0001110000110100", 653 => "1001101010111110", 654 => "1100101101001011", 655 => "1000001110011000", 656 => "0101010111111011", 657 => "1010011010110110", 658 => "1011111011111000", 659 => "1011110111001101", 660 => "1101011101000111", 661 => "0011110000110000", 662 => "1110010001000100", 663 => "0110011000010000", 664 => "0011101101000011", 665 => "0011000000010110", 666 => "0010000001011010", 667 => "0111101010010000", 668 => "1100101011101001", 669 => "0001110110011010", 670 => "1010100011100011", 671 => "1101011001000010", 672 => "1001010010011101", 673 => "1101110111010111", 674 => "1001011010100010", 675 => "1010110100010001", 676 => "1111101110001100", 677 => "0110001110100111", 678 => "0101110101010000", 679 => "1001011100001111", 680 => "0110010101101011", 681 => "0000100101000011", 682 => "0100101111110010", 683 => "0111100000011000", 684 => "1011111101101100", 685 => "1110100010000111", 686 => "0100101100011101", 687 => "1000010010010111", 688 => "1101000001101011", 689 => "1001110100101010", 690 => "1100011101110011", 691 => "1100011110001101", 692 => "0101000000000001", 693 => "1110000010000101", 694 => "0010011010011011", 695 => "0001001011111110", 696 => "0000011101110010", 697 => "1110110101101011", 698 => "1101100101000110", 699 => "0001011111111101", 700 => "1100001100111011", 701 => "0010010001110110", 702 => "0000110100011101", 703 => "1000010000110101", 704 => "0110001011010000", 705 => "1101010000111010", 706 => "0110111110011000", 707 => "0100000100010001", 708 => "0101101111101101", 709 => "1010100110101101", 710 => "0011110110000111", 711 => "0011011111111100", 712 => "0110000001011101", 713 => "1010101111101011", 714 => "1010011001000010", 715 => "1100000110011110", 716 => "1101011011101001", 717 => "0000101111011001", 718 => "1010011100100101", 719 => "0011110001100101", 720 => "1100010101111010", 721 => "1110110011111111", 722 => "1100101000101001", 723 => "1010111101011000", 724 => "0011000001111010", 725 => "0110010001010010", 726 => "1110010010101000", 727 => "1111100011010010", 728 => "0011111111001000", 729 => "1011101111100010", 730 => "0000010101000101", 731 => "0101100111110110", 732 => "0001111000100110", 733 => "0100001111001111", 734 => "0100000100001011", 735 => "0111110011011001", 736 => "0101011011001111", 737 => "1111101110011101", 738 => "0011101000000001", 739 => "1000001110010010", 740 => "0100001010010110", 741 => "1000011011111110", 742 => "1100001111010110", 743 => "0001100110010101", 744 => "1010101000001101", 745 => "1000101110110011", 746 => "0101001100100100", 747 => "0110010011001010", 748 => "1010000100100110", 749 => "0000010010011000", 750 => "0001100111010001", 751 => "1100001111011110", 752 => "0001110100110101", 753 => "1011110011010010", 754 => "0010010100101000", 755 => "1000100101010000", 756 => "1001110000110001", 757 => "1101010011101001", 758 => "0000101011010011", 759 => "0111001110110010", 760 => "0100100101111101", 761 => "1001100000011100", 762 => "0000110110000001", 763 => "0110100001101001", 764 => "1111011001001111", 765 => "0001100011100000", 766 => "1111000011111011", 767 => "0011001001110010", 768 => "0000100000110101", 769 => "1001111000110001", 770 => "1101111010001110", 771 => "1111000010101101", 772 => "1101101101110011", 773 => "0110011000001110", 774 => "1110001011110101", 775 => "1010010110101000", 776 => "0010101011101111", 777 => "1000100100010001", 778 => "1001011100001100", 779 => "1111010111101000", 780 => "0001010001111010", 781 => "1010100111100111", 782 => "1110010101101011", 783 => "1000001001111010", 784 => "1101111010100010", 785 => "1110111000001101", 786 => "1011111100011100", 787 => "0001001110011101", 788 => "1010111010001010", 789 => "0100001001110101", 790 => "0111111110001100", 791 => "0000011100000011", 792 => "0101101011100000", 793 => "0110011011011111", 794 => "1101010101111101", 795 => "1011100001100100", 796 => "1010100111011101", 797 => "0100001111011000", 798 => "1110000000101110", 799 => "0111000101010100", 800 => "1101000001001001", 801 => "0001111101000100", 802 => "1010001001000110", 803 => "0110110000011010", 804 => "0010111001111010", 805 => "0011101000100111", 806 => "1000101000110101", 807 => "1100110100011111", 808 => "1111110111011110", 809 => "0010110101010010", 810 => "0101011101000001", 811 => "0001110011101010", 812 => "1100000011010010", 813 => "0000010001110000", 814 => "1110111101010011", 815 => "1000101101001011", 816 => "0100100110011101", 817 => "1111011111110101", 818 => "0000000101110011", 819 => "0101100101101000", 820 => "1111001011100100", 821 => "0101101100011000", 822 => "1010100010011011", 823 => "0001000100011011", 824 => "0010011110110011", 825 => "1001111010101011", 826 => "0011101001101111", 827 => "1001111110000101", 828 => "0101101111101010", 829 => "0110010101000111", 830 => "0001111000010111", 831 => "1001110000001101", 832 => "1101010111000111", 833 => "0101111100010010", 834 => "1001111000000011", 835 => "0000001011101011", 836 => "1101011100100110", 837 => "1110011001011101", 838 => "0000001110001011", 839 => "1101111000011001", 840 => "0100000001000001", 841 => "1011110100100110", 842 => "0110011001111111", 843 => "1001010111111111", 844 => "1001011101110001", 845 => "0100000000100110", 846 => "0000010110111010", 847 => "1110110000010001", 848 => "1000101111000000", 849 => "1000111001011001", 850 => "1100111100011100", 851 => "1010100010100101", 852 => "0000100001010010", 853 => "1101010100011111", 854 => "0100001110100011", 855 => "1101100000011100", 856 => "1110011010000101", 857 => "0101000001010010", 858 => "0100110001001010", 859 => "1111111011100101", 860 => "0111110101010011", 861 => "0010000010101111", 862 => "1111010011010111", 863 => "1011110100110000", 864 => "0100001000010000", 865 => "1010101010101001", 866 => "0011000111111111", 867 => "0001000011001100", 868 => "1100100011010110", 869 => "1001111000110110", 870 => "1000110000001011", 871 => "1010001011001000", 872 => "0010101100111001", 873 => "0000100000110000", 874 => "0100101110101100", 875 => "1011010110110100", 876 => "0111110001010110", 877 => "0001000110101011", 878 => "1101011000010100", 879 => "1101101110101111", 880 => "0010100110000110", 881 => "1110110111001110", 882 => "1101100100101000", 883 => "1001110110111000", 884 => "1010011101110001", 885 => "0001011001000010", 886 => "0111001011001000", 887 => "0111011111110100", 888 => "0011111101011111", 889 => "0100011100000111", 890 => "1011111011010110", 891 => "0010111011111110", 892 => "1001100011010000", 893 => "0010111001001101", 894 => "1000010010100101", 895 => "0101010011000000", 896 => "0100100111110011", 897 => "0111100001110001", 898 => "1000110001011111", 899 => "0011101001000101", 900 => "0010011100111101", 901 => "1010100110100111", 902 => "1111010000000100", 903 => "0011000011001010", 904 => "0111011111101111", 905 => "1100101010101001", 906 => "1100101111010111", 907 => "0110100010100001", 908 => "1100110010100110", 909 => "0110110010011010", 910 => "0111010111001001", 911 => "0010011101000011", 912 => "0111000000001110", 913 => "1010100111010010", 914 => "1100100001000111", 915 => "0000110011001000", 916 => "0000111100111000", 917 => "1010100111011010", 918 => "1011000000000110", 919 => "0110111010011000", 920 => "0111011001011000", 921 => "1010110110000110", 922 => "0010100000001111", 923 => "0110000011010110", 924 => "1000110010001011", 925 => "1111101001111010", 926 => "1100000001000100", 927 => "0010100110001110", 928 => "1011111011000111", 929 => "0011011011101110", 930 => "1110001001000110", 931 => "1001111100101010", 932 => "0010000010101000", 933 => "1100100000000001", 934 => "1001100101100100", 935 => "1110010010010001", 936 => "0100100110010010", 937 => "0001011011001111", 938 => "0100111011010001", 939 => "1001110110001011", 940 => "0100010110101100", 941 => "1000110110111111", 942 => "0100000111001011", 943 => "1000111110000011", 944 => "1011111001110001", 945 => "1001001101011100", 946 => "0000000111101001", 947 => "0101110100011011", 948 => "0111100010110111", 949 => "0010010110101101", 950 => "1101111000101001", 951 => "1100000001101001", 952 => "0011000011111010", 953 => "1010010001010101", 954 => "0111010001001010", 955 => "1000000000010111", 956 => "0101000010010111", 957 => "1101101001011111", 958 => "1111011001011011", 959 => "1100100101110100", 960 => "1101100001011101", 961 => "0100011010000110", 962 => "0100010011010011", 963 => "0101101100100100", 964 => "0000001101011111", 965 => "0010010011011011", 966 => "0011111001000111", 967 => "0000101000110100", 968 => "1001000000100001", 969 => "1100100101101100", 970 => "0001011100000110", 971 => "0000000011111110", 972 => "1111001011110100", 973 => "0101110000011100", 974 => "0010101010100010", 975 => "1001110000101101", 976 => "1100110100011000", 977 => "1011101000100000", 978 => "0010110001111000", 979 => "1111110110111100", 980 => "1101010110110001", 981 => "0100110001101110", 982 => "1000111110011101", 983 => "1001000111110000", 984 => "0001101101100111", 985 => "0111001000001100", 986 => "1101000011100011", 987 => "0101100001011111", 988 => "1111100100011011", 989 => "1101111001110100", 990 => "1010111001010011", 991 => "0100011011101110", 992 => "1110010110010101", 993 => "0110011011011100", 994 => "0000101111011000", 995 => "0100110001010111", 996 => "0110111000010100", 997 => "1101101111000011", 998 => "1001101001111100", 999 => "0110000010010001", 1000 => "1100010010010011", 1001 => "1000000000011010", 1002 => "0111001001001100", 1003 => "1001010000000111", 1004 => "1100010101111001", 1005 => "1011100011010011", 1006 => "0011110101001101", 1007 => "1001110010111111", 1008 => "1000010100011111", 1009 => "1000001111111000", 1010 => "1101001110010111", 1011 => "1011000001101001", 1012 => "1111010110101111", 1013 => "1111110111001010", 1014 => "0101111101001101", 1015 => "0000111100101101", 1016 => "0111111111000011", 1017 => "0100000110110000", 1018 => "0001010000101001", 1019 => "1011100100000100", 1020 => "0011110011110101", 1021 => "0110101100011111", 1022 => "1010111111101010", 1023 => "1110010101110001", 1024 => "0110100111011010", 1025 => "0101100000111110", 1026 => "1000110111101101", 1027 => "1110000100011100", 1028 => "0001110010100111", 1029 => "1010111101111000", 1030 => "1101010011001101", 1031 => "0111100000110101", 1032 => "1110100010001110", 1033 => "0100100010011000", 1034 => "1110110100100001", 1035 => "1011011100110000", 1036 => "1111100001011101", 1037 => "0101111011011101", 1038 => "1010000011100110", 1039 => "0100101101001011", 1040 => "1111100011010010", 1041 => "0010000011101010", 1042 => "1010100000000000", 1043 => "1100000001110100", 1044 => "1101001111011010", 1045 => "0100111100011100", 1046 => "1001011101011111", 1047 => "1101011101010011", 1048 => "1010010011101111", 1049 => "0000011000010010", 1050 => "0001011001000100", 1051 => "0010100010101000", 1052 => "0010101011010110", 1053 => "1011110110001011", 1054 => "0111110001110111", 1055 => "0001011000001010", 1056 => "0000111100011001", 1057 => "1011000100000100", 1058 => "1000001110111100", 1059 => "0111000011110001", 1060 => "0011000001001100", 1061 => "0011010011101100", 1062 => "1110111110111100", 1063 => "1111001011001010", 1064 => "0001100100000110", 1065 => "0100001011011111", 1066 => "0001000000100111", 1067 => "0011000010010001", 1068 => "1001011011111101", 1069 => "0011010111011010", 1070 => "0011010011001111", 1071 => "0100100111000111", 1072 => "0101101100101010", 1073 => "1000000110010111", 1074 => "0111010100001010", 1075 => "1011110010010011", 1076 => "1110001010010100", 1077 => "1001001000000111", 1078 => "1101010001100011", 1079 => "0000111010010100", 1080 => "0011010111010010", 1081 => "1000011000011101", 1082 => "0111101110101000", 1083 => "0100001010000110", 1084 => "0100011001011000", 1085 => "0101000101111110", 1086 => "1011100100111000", 1087 => "1110111101111001", 1088 => "0001100010101000", 1089 => "1110111001001010", 1090 => "0011101011101011", 1091 => "1100100100100110", 1092 => "1010011111000100", 1093 => "1111011111010100", 1094 => "1011001100001110", 1095 => "0110000101000101", 1096 => "0010000010001001", 1097 => "1000111100111000", 1098 => "1100010100001010", 1099 => "0010001001001010", 1100 => "1010101101111111", 1101 => "1110100101011100", 1102 => "0101000101001101", 1103 => "1110010001010011", 1104 => "1111110100101110", 1105 => "1111100000100011", 1106 => "1011111001001110", 1107 => "1011001011010001", 1108 => "0000001111010100", 1109 => "0110100101001101", 1110 => "1100001001100110", 1111 => "1000101000111001", 1112 => "1000110101011010", 1113 => "1000011001110010", 1114 => "1000111110101000", 1115 => "0000110100010000", 1116 => "1011101101111100", 1117 => "0000110000111010", 1118 => "1010111110110001", 1119 => "0101001010101111", 1120 => "1111100000100010", 1121 => "0111100000111100", 1122 => "1011111011101010", 1123 => "1101011111001010", 1124 => "1011001011100100", 1125 => "1011000110011010", 1126 => "1001000010011001", 1127 => "1010110110011100", 1128 => "0111100010110100", 1129 => "0110010000100000", 1130 => "1111010000011111", 1131 => "0011011111011111", 1132 => "0011010011000101", 1133 => "0010100100001000", 1134 => "0110001000000100", 1135 => "0001010011111110", 1136 => "1100010111000011", 1137 => "0111011110110000", 1138 => "0001110010100110", 1139 => "1000001001110101", 1140 => "1101000110101010", 1141 => "0010001111101010", 1142 => "0000111100101011", 1143 => "1101010000010111", 1144 => "1001001101011011", 1145 => "1110011100110100", 1146 => "1000011101111101", 1147 => "0111100011001101", 1148 => "1110110111101011", 1149 => "1010101011111001", 1150 => "0010110001110100", 1151 => "1100001100111110", 1152 => "0101001010011011", 1153 => "0011000111011101", 1154 => "0000011011001001", 1155 => "0010010100010001", 1156 => "1101010010010010", 1157 => "1111111011011101", 1158 => "1101101000011001", 1159 => "1101101101001111", 1160 => "0000100111001100", 1161 => "0110010101011111", 1162 => "0110101110001100", 1163 => "0111111110001011", 1164 => "0010010110010001", 1165 => "0001001101001101", 1166 => "0110001100100011", 1167 => "0001111010111101", 1168 => "0001110101101101", 1169 => "0000100111001000", 1170 => "1111000010111011", 1171 => "1111100111101100", 1172 => "0010101111001011", 1173 => "1101010000110110", 1174 => "0010110000100000", 1175 => "1110011101010000", 1176 => "1000111011011000", 1177 => "1100110010001101", 1178 => "0001100111111110", 1179 => "0011111010110101", 1180 => "0101111010000111", 1181 => "1111010011001010", 1182 => "0010110001101001", 1183 => "0000000101111100", 1184 => "1011110110110001", 1185 => "0110000011001101", 1186 => "0011011110110010", 1187 => "0011110001110111", 1188 => "1010100000100001", 1189 => "1010101100101001", 1190 => "0101011111010101", 1191 => "0111000011000011", 1192 => "0010100101110000", 1193 => "0111011011111111", 1194 => "0010100110101111", 1195 => "1011001111101101", 1196 => "0001011000101011", 1197 => "0010010010001101", 1198 => "0010010101011011", 1199 => "1100000011111100", 1200 => "1000101101011111", 1201 => "1010101001101011", 1202 => "1101100111101011", 1203 => "0011101010011111", 1204 => "1000100110011001", 1205 => "0101001110010010", 1206 => "0100001111000101", 1207 => "0111010110011000", 1208 => "1010111111101010", 1209 => "1110100001101000", 1210 => "1101000011011000", 1211 => "1010011101000000", 1212 => "1010110110000100", 1213 => "0001111000110011", 1214 => "1001001110100101", 1215 => "1111101011001001", 1216 => "1000111010111110", 1217 => "0111001001101001", 1218 => "0110111010001010", 1219 => "0101110000101001", 1220 => "1100100010111001", 1221 => "1011000100000001", 1222 => "1100111000011010", 1223 => "1111101110110011", 1224 => "0000001110110010", 1225 => "1001110111111110", 1226 => "0101011000010101", 1227 => "0101000111010001", 1228 => "1111100111000001", 1229 => "1110010111001001", 1230 => "0011111010000111", 1231 => "1101110000100011", 1232 => "1000010010110111", 1233 => "0100000011101000", 1234 => "0001000010110100", 1235 => "0101000101111001", 1236 => "0110010101111011", 1237 => "1010000001000101", 1238 => "1111011000111100", 1239 => "0011111000111111", 1240 => "0011100111110011", 1241 => "0001010100101000", 1242 => "0100100101110011", 1243 => "1101000011110101", 1244 => "0110100011011111", 1245 => "1000111010001001", 1246 => "0110000101001001", 1247 => "0110000000100000", 1248 => "0110010000010100", 1249 => "0100000011110000", 1250 => "1000110110000000", 1251 => "1001101000001010", 1252 => "0101101010111110", 1253 => "1010010101000010", 1254 => "0100110001011110", 1255 => "1011001100010100", 1256 => "1100101111100001", 1257 => "1011110011011000", 1258 => "0011001000101101", 1259 => "1110111001100100", 1260 => "0010100001110100", 1261 => "1111101001000100", 1262 => "0111101001111100", 1263 => "1111001100111110", 1264 => "0011110001110100", 1265 => "1111001000011100", 1266 => "0010100100011001", 1267 => "1000001101001001", 1268 => "0110101001011110", 1269 => "0011011011111110", 1270 => "0000011000110000", 1271 => "1000110001110011", 1272 => "1100100101111010", 1273 => "0111110100010110", 1274 => "1001100010011001", 1275 => "1000100110001010", 1276 => "0010111011011001", 1277 => "1001100000001111", 1278 => "0011111001010010", 1279 => "1100001010010111", 1280 => "1110101100001000", 1281 => "1011010000111111", 1282 => "1100011100010001", 1283 => "1101000011110010", 1284 => "0010000110011010", 1285 => "0110110101000001", 1286 => "0011100101100000", 1287 => "1001110000111111", 1288 => "1010111000110000", 1289 => "1001101001111010", 1290 => "0000011111110001", 1291 => "1001010110110101", 1292 => "1000110111001011", 1293 => "0000001010010101", 1294 => "0011110101111000", 1295 => "1110001101011000", 1296 => "1110111111011100", 1297 => "1100111110111100", 1298 => "1000101111110101", 1299 => "0001100110101000", 1300 => "0111000111001101", 1301 => "1010011100101110", 1302 => "1001101000111110", 1303 => "0101111110111110", 1304 => "0011110111000001", 1305 => "0100100011110100", 1306 => "0100011111000110", 1307 => "1100011001101010", 1308 => "0000111110010101", 1309 => "1100100000101101", 1310 => "0101001001001001", 1311 => "0111011100010100", 1312 => "1111111111111001", 1313 => "0101111110001000", 1314 => "0001001101100010", 1315 => "1000100110101100", 1316 => "1111000111011010", 1317 => "0101001000101001", 1318 => "0011010011110101", 1319 => "1010011011000000", 1320 => "0011110011100101", 1321 => "0001100001101101", 1322 => "0000100100000101", 1323 => "1110101000100010", 1324 => "1010110010001010", 1325 => "1111001100000000", 1326 => "1110011011010110", 1327 => "0000101110001000", 1328 => "0011111111100101", 1329 => "1001000010000101", 1330 => "0010110010011110", 1331 => "1110001011011101", 1332 => "0111100001101100", 1333 => "0110101010010000", 1334 => "0000001101101110", 1335 => "0100111110110010", 1336 => "1010000101000100", 1337 => "1001110010111011", 1338 => "0011010000110001", 1339 => "0001100101110011", 1340 => "0111111101010101", 1341 => "0010001110011110", 1342 => "1001110110010111", 1343 => "1000111011111000", 1344 => "1111011011001100", 1345 => "0000110101101001", 1346 => "1110011110111110", 1347 => "0000001111010000", 1348 => "0110010010101101", 1349 => "0011001001101000", 1350 => "0100110100011110", 1351 => "0100000101100100", 1352 => "1001011101111100", 1353 => "1001000011110100", 1354 => "1101111011011000", 1355 => "0111010010110111", 1356 => "0100101111000001", 1357 => "0010110110000100", 1358 => "1110100010110100", 1359 => "0100101111110110", 1360 => "1000010111010101", 1361 => "0111000101001101", 1362 => "0100011011101101", 1363 => "0110110100001101", 1364 => "0101101010110100", 1365 => "1110110100110111", 1366 => "0110111001000110", 1367 => "1011110100100001", 1368 => "0100111101101101", 1369 => "0001010100101100", 1370 => "0100111001001001", 1371 => "1110010001111001", 1372 => "0010101100110010", 1373 => "1011011101011101", 1374 => "0111010001111100", 1375 => "0000111001011101", 1376 => "1010100110000111", 1377 => "1100100110111010", 1378 => "1010011101001110", 1379 => "1011000010000000", 1380 => "0101100110111010", 1381 => "0100000000011011", 1382 => "0001010001111001", 1383 => "0111010011110110", 1384 => "1100110111011111", 1385 => "0011011100001100", 1386 => "1000100111000000", 1387 => "0010110100111001", 1388 => "0101000101000101", 1389 => "1100100011101000", 1390 => "1011111111111010", 1391 => "0100010101011001", 1392 => "0110000100001101", 1393 => "1101000010100110", 1394 => "0001111111001100", 1395 => "0010101101101000", 1396 => "1110100001101101", 1397 => "0000001000101000", 1398 => "0011100100110011", 1399 => "0111101001010110", 1400 => "1101110010110000", 1401 => "0010111011010001", 1402 => "0101101000001100", 1403 => "0010110101110110", 1404 => "1100011110111011", 1405 => "0100011101111100", 1406 => "1001110111101111", 1407 => "1011110101010101", 1408 => "1011101010101010", 1409 => "0111010100001100", 1410 => "0101011111100111", 1411 => "1110101011011110", 1412 => "1001010111000110", 1413 => "1110111010101001", 1414 => "1011000000101011", 1415 => "0001001001111000", 1416 => "1000101010100101", 1417 => "0001010101001001", 1418 => "1111010011100101", 1419 => "0011101111111100", 1420 => "1100001011110010", 1421 => "1110010011011110", 1422 => "1011100100101010", 1423 => "1111011001111010", 1424 => "1011111111010011", 1425 => "0000111001011001", 1426 => "0000001001110100", 1427 => "1111000010000111", 1428 => "0110000111000010", 1429 => "1100100101111100", 1430 => "0100001011011101", 1431 => "0011111111000000", 1432 => "0111010101000000", 1433 => "1100011111001010", 1434 => "0111000010010101", 1435 => "1011000011001110", 1436 => "0011101110101100", 1437 => "1000000011000101", 1438 => "1110010001101110", 1439 => "1000010001111100", 1440 => "0000111100101101", 1441 => "1000010001011001", 1442 => "0000010100010010", 1443 => "0100110101110001", 1444 => "0001001101110001", 1445 => "1110110110111011", 1446 => "0000010110011111", 1447 => "0010110110111001", 1448 => "1111001011101000", 1449 => "0000110001011111", 1450 => "0111100010111010", 1451 => "0000111101100101", 1452 => "1110101100000100", 1453 => "1011000111010101", 1454 => "1100111100011011", 1455 => "1011110101001011", 1456 => "1110111000000001", 1457 => "1100010011000101", 1458 => "1001101011000100", 1459 => "1100001110010111", 1460 => "1000110001110001", 1461 => "0111001010011011", 1462 => "0010110001000010", 1463 => "0110100010011111", 1464 => "0101110010011110", 1465 => "1000111101000001", 1466 => "0111110011010011", 1467 => "0110100111101001", 1468 => "0001110111010101", 1469 => "1001000100010101", 1470 => "0000011111011100", 1471 => "0000001010010001", 1472 => "0101011101001100", 1473 => "1001101000011001", 1474 => "0110010110111001", 1475 => "1001010011111000", 1476 => "1110000111100101", 1477 => "1000111010110010", 1478 => "1111100110101111", 1479 => "1111110011011101", 1480 => "0000111100100000", 1481 => "0110111001101001", 1482 => "1010100011101110", 1483 => "0111111010000111", 1484 => "1100100111010101", 1485 => "0111010110011101", 1486 => "1111100110000111", 1487 => "1000110101101010", 1488 => "1011111101001001", 1489 => "0001100100001101", 1490 => "1100001110011110", 1491 => "1000000011010111", 1492 => "1101000000011011", 1493 => "1011101111110100", 1494 => "1100010101010100", 1495 => "1111100011100110", 1496 => "0010101001010110", 1497 => "0111111000100100", 1498 => "0100010100011110", 1499 => "0110001001010010", 1500 => "0110100110010011", 1501 => "1100001110011100", 1502 => "1110100000101010", 1503 => "0101011110011000", 1504 => "0110110000011000", 1505 => "1000001100100111", 1506 => "1100111010111000", 1507 => "0100000000001101", 1508 => "0011100100011001", 1509 => "0010110110010001", 1510 => "1111000111111111", 1511 => "1011001011110111", 1512 => "1001000110010101", 1513 => "1111101101110011", 1514 => "0011010011001010", 1515 => "1010000110010010", 1516 => "0001110100100101", 1517 => "0111101111011000", 1518 => "1101011100000000", 1519 => "0010000101011010", 1520 => "0010100111110100", 1521 => "0111111001111000", 1522 => "0111100111010101", 1523 => "1011101001101100", 1524 => "0101100111010001", 1525 => "0100001100101110", 1526 => "1010110101011010", 1527 => "1010001111011000", 1528 => "1001001010010000", 1529 => "0011111111010101", 1530 => "0100100010111010", 1531 => "0100110010110101", 1532 => "1100110100010111", 1533 => "1110000110011111", 1534 => "0000110100010100", 1535 => "1110001110001010", 1536 => "0100010100010111", 1537 => "0000110100110100", 1538 => "1111100010111111", 1539 => "0100010011010100", 1540 => "1001110100000010", 1541 => "0000111001010111", 1542 => "0110100111000010", 1543 => "1101111011000100", 1544 => "1000111111101011", 1545 => "1101100101101101", 1546 => "1001111010101000", 1547 => "0101010111101100", 1548 => "0111010010101110", 1549 => "1111010110001000", 1550 => "1111000010000100", 1551 => "1000111001010001", 1552 => "0001010111010111", 1553 => "0000101101110010", 1554 => "1110000000101001", 1555 => "0100001110101000", 1556 => "0010101001000101", 1557 => "0101000011011111", 1558 => "0110001101010000", 1559 => "0010101100000000", 1560 => "0001001000100011", 1561 => "1110011011011110", 1562 => "1011101000111001", 1563 => "0011110111011111", 1564 => "0010000111001000", 1565 => "0000111011111110", 1566 => "1000010110011010", 1567 => "1001110011010011", 1568 => "1101001011101101", 1569 => "1000000111100010", 1570 => "0011001111011101", 1571 => "1111010000011100", 1572 => "1101001001101001", 1573 => "1110100101001100", 1574 => "1011111000011010", 1575 => "1010101110111101", 1576 => "1011111101101101", 1577 => "1011111111000100", 1578 => "1000101101000110", 1579 => "1010001110000100", 1580 => "1110111100101100", 1581 => "1010010110111111", 1582 => "0001100100100000", 1583 => "0011110010011000", 1584 => "1111000001001111", 1585 => "1110010110101000", 1586 => "0001010110010011", 1587 => "1000000000001001", 1588 => "0001110111010010", 1589 => "1100001100100011", 1590 => "0110110011010001", 1591 => "0111000011000000", 1592 => "1110101101010011", 1593 => "1011101001001001", 1594 => "0111100100001010", 1595 => "0010000101010101", 1596 => "0000001100100110", 1597 => "1001000011110010", 1598 => "1100011011100001", 1599 => "0001010110010011", 1600 => "1100111111100001", 1601 => "1101101001001100", 1602 => "0100001110101101", 1603 => "0001110111100011", 1604 => "1111000100100100", 1605 => "0110011011111010", 1606 => "0011001110101010", 1607 => "1100001010010001", 1608 => "0101110000000110", 1609 => "1100000010000110", 1610 => "1100000000011001", 1611 => "0101111010110000", 1612 => "1000000101011101", 1613 => "0100101100000101", 1614 => "0011111000010110", 1615 => "0000011011010110", 1616 => "1010111111110010", 1617 => "0001100000001001", 1618 => "0110110100000100", 1619 => "1101001110001100", 1620 => "0101011101100000", 1621 => "1110001010100100", 1622 => "1100001100110110", 1623 => "1110000101010100", 1624 => "0011111100111011", 1625 => "0110100000000010", 1626 => "0010010101010101", 1627 => "0000000001010110", 1628 => "1100010100111101", 1629 => "1011100110111000", 1630 => "1110010010011101", 1631 => "0011101001101001", 1632 => "0000110101001101", 1633 => "1110110010111111", 1634 => "0010011010110101", 1635 => "0101110001101010", 1636 => "1000000110100110", 1637 => "1110101110111011", 1638 => "1001001111010100", 1639 => "0111101000110100", 1640 => "1001000001101101", 1641 => "0110111001010111", 1642 => "1101001100101001", 1643 => "1110100100100000", 1644 => "1011011111101101", 1645 => "0001001001100101", 1646 => "1100001110111001", 1647 => "0110111001111011", 1648 => "0011011100001011", 1649 => "0111100110110011", 1650 => "1011111001111000", 1651 => "0010010000000000", 1652 => "1100111010111100", 1653 => "1111100011010100", 1654 => "0100101111100111", 1655 => "0011110000001001", 1656 => "0100111101000100", 1657 => "0011000110101111", 1658 => "0000001111011100", 1659 => "1010110110101011", 1660 => "1101010110110110", 1661 => "1111001000011111", 1662 => "0111100001011100", 1663 => "0101001100110001", 1664 => "1011001001100111", 1665 => "0101111110111011", 1666 => "1111100111101101", 1667 => "0010010011000010", 1668 => "0100100001111110", 1669 => "0010011110111001", 1670 => "0110100011110100", 1671 => "1001101011101110", 1672 => "0011110101011111", 1673 => "0001100001001000", 1674 => "0101101001000000", 1675 => "1010011110011100", 1676 => "0011110000001101", 1677 => "0100010110101011", 1678 => "1000011000111000", 1679 => "1011010000111010", 1680 => "1000111110100001", 1681 => "1101001000101001", 1682 => "1100101011100110", 1683 => "1010000011001100", 1684 => "0110110010011110", 1685 => "0101111000101110", 1686 => "1100011101111011", 1687 => "1111000100010111", 1688 => "0101000111000011", 1689 => "0100100011110011", 1690 => "1101010101101011", 1691 => "0001000100111010", 1692 => "1010011011001001", 1693 => "0001111100010010", 1694 => "1101101101111110", 1695 => "0001111011101111", 1696 => "1000101011111110", 1697 => "1001001100011111", 1698 => "1110110101000010", 1699 => "1101001101111000", 1700 => "0010110000100011", 1701 => "0001000010101000", 1702 => "1101001010101111", 1703 => "1111001110101010", 1704 => "1101110100100011", 1705 => "0101101111111100", 1706 => "1011010000101011", 1707 => "1101111110011110", 1708 => "1001010000000011", 1709 => "0001111111001011", 1710 => "1010001100000110", 1711 => "0111101011001011", 1712 => "0011000111000011", 1713 => "0111001010010011", 1714 => "1001110101000100", 1715 => "1110000010010111", 1716 => "1001000011101010", 1717 => "1000100001111101", 1718 => "0101000100010000", 1719 => "0011010011000000", 1720 => "0101110101000101", 1721 => "1110101000101110", 1722 => "0111010110001000", 1723 => "0100111111111001", 1724 => "0110100000010111", 1725 => "1110110010100000", 1726 => "0000011001110000", 1727 => "1111000010101011", 1728 => "0101110110000011", 1729 => "0010011000011001", 1730 => "1001010000111101", 1731 => "0011110101010111", 1732 => "0111111110101110", 1733 => "0111101110011111", 1734 => "1111010111011110", 1735 => "0100100110101001", 1736 => "0110110000100001", 1737 => "0010111000000010", 1738 => "1001001000101100", 1739 => "1010110011000000", 1740 => "1001100011001110", 1741 => "0110101110110001", 1742 => "0110110110101101", 1743 => "0011100100101101", 1744 => "1001100011111111", 1745 => "0011000010011000", 1746 => "1001110000100001", 1747 => "0110011000001111", 1748 => "1111011100100101", 1749 => "0110010101000011", 1750 => "1111010001111000", 1751 => "1101110010110010", 1752 => "0011010111011110", 1753 => "1100100011000010", 1754 => "1101000000100000", 1755 => "1000111101101101", 1756 => "0010000001111100", 1757 => "0000110101110110", 1758 => "1011000011010100", 1759 => "0010110101111111", 1760 => "0101010000011000", 1761 => "0101010100110110", 1762 => "1110101111100101", 1763 => "1000011100010110", 1764 => "0000100111110011", 1765 => "1111000001101011", 1766 => "1110101000111011", 1767 => "0110010000100011", 1768 => "1101011000001000", 1769 => "1011111110011100", 1770 => "0010110001001110", 1771 => "0111010111111101", 1772 => "1110011100100011", 1773 => "1001111010000011", 1774 => "0111000111100110", 1775 => "1011110010001111", 1776 => "0000001000001100", 1777 => "0000101110011011", 1778 => "0001101000001010", 1779 => "0010001100110100", 1780 => "1001011110000000", 1781 => "1000000101110011", 1782 => "1111010100100011", 1783 => "1111011111101011", 1784 => "1011000110010000", 1785 => "0010111101101001", 1786 => "1100111000101110", 1787 => "0000010010001001", 1788 => "1011000011111000", 1789 => "0111101011000100", 1790 => "1111110110111101", 1791 => "0001001110010011", 1792 => "0001000011010100", 1793 => "1010110010110111", 1794 => "1000000101001001", 1795 => "0000000110001001", 1796 => "0011010111001110", 1797 => "1001001110110111", 1798 => "1010110001010101", 1799 => "1110001011001100", 1800 => "0001111100010011", 1801 => "0100110011100111", 1802 => "0111001000101110", 1803 => "1111011110101011", 1804 => "1001110010001101", 1805 => "1110010010111000", 1806 => "0010001101111111", 1807 => "1111010000000111", 1808 => "0100110101101000", 1809 => "0010111011011101", 1810 => "0000011110110101", 1811 => "1000111010110111", 1812 => "0101110111011011", 1813 => "0001011011000110", 1814 => "0101100000001101", 1815 => "1000001001001001", 1816 => "1101100100111101", 1817 => "0000101101111110", 1818 => "0101100100010110", 1819 => "1011011111010101", 1820 => "1010000000100111", 1821 => "0010010010111000", 1822 => "0100111010001010", 1823 => "0000000011000011", 1824 => "1011100001100111", 1825 => "0000101011110101", 1826 => "0010101111010100", 1827 => "0010010000100010", 1828 => "0011111110100000", 1829 => "0100000100100110", 1830 => "0000110111001001", 1831 => "1001111001011111", 1832 => "0110111000011110", 1833 => "0100010110001101", 1834 => "1101110011001000", 1835 => "0101011111010111", 1836 => "0011100111101111", 1837 => "1010110110010101", 1838 => "1100111010111001", 1839 => "1110101111001111", 1840 => "0011100010101111", 1841 => "0110000111110011", 1842 => "1110111100011000", 1843 => "0110110001010001", 1844 => "0111011110110101", 1845 => "0001011011001110", 1846 => "0011010111010100", 1847 => "0101000011101011", 1848 => "0010101100100001", 1849 => "1001010001000111", 1850 => "1110001101110111", 1851 => "1011110011011100", 1852 => "0011001101100000", 1853 => "0001111000001001", 1854 => "0011010010101000", 1855 => "0110001110010111", 1856 => "0011011111001000", 1857 => "0010010100101001", 1858 => "1100011001101011", 1859 => "0010001001001010", 1860 => "1110100010101001", 1861 => "1000010111010000", 1862 => "1001011110100111", 1863 => "1111100110001110", 1864 => "0101010101101000", 1865 => "0111101011010100", 1866 => "0001000101001111", 1867 => "0100111011000010", 1868 => "0000000011011001", 1869 => "0100001011101010", 1870 => "0000011001101101", 1871 => "1101101001100110", 1872 => "1011000011001110", 1873 => "1110100100010101", 1874 => "0111110010000011", 1875 => "0100110001001110", 1876 => "1101010000001000", 1877 => "1000010001010101", 1878 => "0011111110000010", 1879 => "0010100000111001", 1880 => "1011001001101110", 1881 => "0101111001011011", 1882 => "1011001111100101", 1883 => "1110100100101100", 1884 => "0011001011010011", 1885 => "1100101101110100", 1886 => "1100110001111101", 1887 => "1000110100100000", 1888 => "1101001000010111", 1889 => "1011001010010111", 1890 => "0101111100111101", 1891 => "0100110011111100", 1892 => "1110101100101001", 1893 => "1100100010100100", 1894 => "0001000010010101", 1895 => "0001101010110111", 1896 => "1101101110000011", 1897 => "0011011001100101", 1898 => "0010001011000100", 1899 => "1000000110111111", 1900 => "0001100101001011", 1901 => "1101100011010110", 1902 => "0100010110010001", 1903 => "1110010011011001", 1904 => "0110111011001101", 1905 => "1010100100001100", 1906 => "1100110101101100", 1907 => "0010101001111011", 1908 => "0111000011101011", 1909 => "0001011101100011", 1910 => "1111001010101000", 1911 => "0111010011011100", 1912 => "1111110110010110", 1913 => "0001100111011110", 1914 => "0001000011010000", 1915 => "0011100010111001", 1916 => "1011001111001110", 1917 => "1011111100100111", 1918 => "0001100011011110", 1919 => "1000111001000101", 1920 => "1101111110000010", 1921 => "0010111001000000", 1922 => "0010110101001110", 1923 => "1111100111100001", 1924 => "1111010100010101", 1925 => "1001101101010001", 1926 => "1111110110111100", 1927 => "0010010100000101", 1928 => "1000010000000011", 1929 => "1110001000011100", 1930 => "0101011110100111", 1931 => "1010111101100011", 1932 => "1111100001010101", 1933 => "0110101110101110", 1934 => "1100001101110011", 1935 => "1111000001101001", 1936 => "1000110101010111", 1937 => "0110111110001101", 1938 => "0110100010000111", 1939 => "0110111000100110", 1940 => "0100010001001100", 1941 => "1101101011110101", 1942 => "1111001101011011", 1943 => "0011000010000110", 1944 => "0001101110001001", 1945 => "1000111110110110", 1946 => "0011110010110101", 1947 => "1001110011110100", 1948 => "0100100001111000", 1949 => "0000110101000010", 1950 => "1111100111101110", 1951 => "0111000010111001", 1952 => "0110001000110001", 1953 => "1110101010111011", 1954 => "0100100111011111", 1955 => "0001100001101000", 1956 => "1001001110110110", 1957 => "1101011110100100", 1958 => "1101111111001001", 1959 => "1100111101100101", 1960 => "1000100110011010", 1961 => "1010100010000101", 1962 => "0010100010000000", 1963 => "0001101011001110", 1964 => "0010001111111011", 1965 => "0100001011100110", 1966 => "0000001011001010", 1967 => "1101011011111100", 1968 => "0100001000101011", 1969 => "0111001101100001", 1970 => "0001011011111101", 1971 => "0110111000110000", 1972 => "0100110101000000", 1973 => "1011100111101111", 1974 => "1011010001010011", 1975 => "1000100110000001", 1976 => "0000001101001000", 1977 => "1010110001000000", 1978 => "1101111101111101", 1979 => "1110110010110101", 1980 => "1001000010011001", 1981 => "1100110000011001", 1982 => "0000100111000110", 1983 => "1001011011001001", 1984 => "1001101011111011", 1985 => "0111011111100000", 1986 => "1000100100000100", 1987 => "0000001010000111", 1988 => "0011100000101000", 1989 => "0001101011101101", 1990 => "0010100011000000", 1991 => "1010001110011000", 1992 => "0010001101110100", 1993 => "0011111011100011", 1994 => "1110100100000101", 1995 => "0111101010101100", 1996 => "0100110101110000", 1997 => "1000100001001001", 1998 => "1111100110101001", 1999 => "0100111010111110", 2000 => "1010110000001001", 2001 => "0000011001100011", 2002 => "1111100100101111", 2003 => "1010001100001011", 2004 => "0101110110010000", 2005 => "1001110000011100", 2006 => "1110001011010100", 2007 => "0100100101010000", 2008 => "1111111001111111", 2009 => "0001011011100011", 2010 => "0100010110000100", 2011 => "1111111001100110", 2012 => "1101000101100010", 2013 => "1000110111110000", 2014 => "1001111001111100", 2015 => "1010111110001001", 2016 => "1000101011110100", 2017 => "0000001001111010", 2018 => "0011010001111000", 2019 => "1111111111111001", 2020 => "1101101100010011", 2021 => "1000100100110001", 2022 => "0001011011000011", 2023 => "0001001011001110", 2024 => "1010000000011010", 2025 => "0101001101101101", 2026 => "1011100110100011", 2027 => "1100100001101000", 2028 => "1111001001010001", 2029 => "0110101001001110", 2030 => "1110001010101000", 2031 => "0011101000100000", 2032 => "1111100110110110", 2033 => "0110000001000111", 2034 => "1001101001001111", 2035 => "0000101011101111", 2036 => "0110110100110010", 2037 => "1001000001011001", 2038 => "1110111001100101", 2039 => "0100010000111111", 2040 => "0111000001100101", 2041 => "1111111100000011", 2042 => "0111000111111010", 2043 => "0110100011000100", 2044 => "0110101010110011", 2045 => "1000101000000011", 2046 => "0010000011010000", 2047 => "0010110001001011", 2048 => "0010010011111101", 2049 => "0111010010001100", 2050 => "0000110011101001", 2051 => "1000011111001000", 2052 => "1100001010000011", 2053 => "0001100010001111", 2054 => "0100000010010110", 2055 => "1010011000101011", 2056 => "0110001101111010", 2057 => "0010001011101010", 2058 => "0001001001101010", 2059 => "0110010110000111", 2060 => "0000010111111011", 2061 => "1110010111011000", 2062 => "1110000100110010", 2063 => "1111110000110111", 2064 => "0001101110101100", 2065 => "1111111011001100", 2066 => "0000011100000000", 2067 => "0110101000111011", 2068 => "1010100000111000", 2069 => "0101101010011111", 2070 => "1111001110101011", 2071 => "1101100010101101", 2072 => "1011011100111010", 2073 => "0000111010100111", 2074 => "0111011110111000", 2075 => "0011000100100010", 2076 => "1110101100000001", 2077 => "1011111000011011", 2078 => "0001011010001111", 2079 => "0010110110101111", 2080 => "1101111010010100", 2081 => "0110001011000100", 2082 => "1111001001110110", 2083 => "0001010111000100", 2084 => "1010001001011011", 2085 => "1000000101110000", 2086 => "0110100010110111", 2087 => "1011010001101111", 2088 => "0110011000111101", 2089 => "0100001010110101", 2090 => "0101001010101001", 2091 => "1011001000011100", 2092 => "0001100010001110", 2093 => "0011011000010110", 2094 => "1010111100100001", 2095 => "1000100011010011", 2096 => "0001111111010101", 2097 => "0001100010011110", 2098 => "1100101110111000", 2099 => "1100001110111111", 2100 => "0110001110011101", 2101 => "0001100110011111", 2102 => "1000011110001110", 2103 => "0011000100110101", 2104 => "1011010110110101", 2105 => "1101111000000110", 2106 => "0101011000011111", 2107 => "0001010111011010", 2108 => "1011101101000001", 2109 => "1011010111100100", 2110 => "1100010111001101", 2111 => "0010011100000000", 2112 => "0101000101100101", 2113 => "0000001000011101", 2114 => "0101110100001111", 2115 => "1010101101010001", 2116 => "1110010000010111", 2117 => "1010001011010101", 2118 => "0000111110100011", 2119 => "0010001111110000", 2120 => "0011111011001010", 2121 => "1100101111101011", 2122 => "1100010010000000", 2123 => "0001010111100000", 2124 => "0011100110000111", 2125 => "0001011011001110", 2126 => "0111110101001101", 2127 => "1100000111110010", 2128 => "0011010100100101", 2129 => "1011001001111101", 2130 => "1100010001100011", 2131 => "1010011100100001", 2132 => "1110101010000000", 2133 => "0101000111011000", 2134 => "1010110010010111", 2135 => "1000110100110110", 2136 => "0100000010000111", 2137 => "0001011011000110", 2138 => "0101100010001110", 2139 => "1101100000100010", 2140 => "1001100000011101", 2141 => "0000110100000101", 2142 => "0010101101011101", 2143 => "0101110001000110", 2144 => "0011000110100110", 2145 => "0110110010000100", 2146 => "1100110011001001", 2147 => "1100101100100100", 2148 => "1100101010001110", 2149 => "0100010101011111", 2150 => "0110011111010100", 2151 => "1011010101111101", 2152 => "0000001111110110", 2153 => "1011010110100101", 2154 => "1011000111011101", 2155 => "0111000010000011", 2156 => "0011001110011001", 2157 => "1011101011011010", 2158 => "0000101111101001", 2159 => "0110111110000100", 2160 => "1010000000010011", 2161 => "1000111111111011", 2162 => "1101000111111001", 2163 => "0010010000111111", 2164 => "1110000101100011", 2165 => "1111100110011000", 2166 => "0001111110100000", 2167 => "1111101011000100", 2168 => "1000000001000111", 2169 => "0111100001011001", 2170 => "0100010100101100", 2171 => "1011000100111110", 2172 => "0100011001111100", 2173 => "1001001001100001", 2174 => "1110100010000011", 2175 => "0111011111001100", 2176 => "1000111100111110", 2177 => "1001010110111111", 2178 => "0011101000001110", 2179 => "0111011000111000", 2180 => "1000101100011100", 2181 => "1000101101101001", 2182 => "1101001110101101", 2183 => "0000100111100000", 2184 => "1110101001110111", 2185 => "1000100101110101", 2186 => "1100001000100101", 2187 => "0110101101001101", 2188 => "0101100100111111", 2189 => "0001011101101000", 2190 => "1100011000000111", 2191 => "0011010110100100", 2192 => "0110011111011100", 2193 => "0111000101001010", 2194 => "0011011101010100", 2195 => "1010001100101011", 2196 => "1101000001100101", 2197 => "1001011001110001", 2198 => "1110011011001101", 2199 => "0101001111110011", 2200 => "0111111111000101", 2201 => "1011110010111011", 2202 => "1110111110101011", 2203 => "1010010111000100", 2204 => "0100001010110111", 2205 => "0010101000001010", 2206 => "0011100110011111", 2207 => "0101000000110100", 2208 => "1001110010010101", 2209 => "0010101011000100", 2210 => "1010011011011000", 2211 => "0001101001101001", 2212 => "1001101011010101", 2213 => "1000101100010110", 2214 => "1000110111101001", 2215 => "0100111111010000", 2216 => "1101000111100110", 2217 => "0101011001010100", 2218 => "0011110001001100", 2219 => "0110110001111011", 2220 => "1000100000110011", 2221 => "1011011101101000", 2222 => "1100100000001001", 2223 => "0100101000010010", 2224 => "1101011101001000", 2225 => "0110111010111101", 2226 => "0111010100011100", 2227 => "1100001001100110", 2228 => "0001110011011001", 2229 => "0000000101101101", 2230 => "1011110100001111", 2231 => "0001010111101111", 2232 => "1010000110010101", 2233 => "1110001100100011", 2234 => "0011110011010000", 2235 => "0111111001100101", 2236 => "0101010011110100", 2237 => "1111111100110000", 2238 => "1110101001010000", 2239 => "1000110011000101", 2240 => "0010010011010110", 2241 => "1110110010001000", 2242 => "1010110100110001", 2243 => "1011000111111101", 2244 => "0001100001010010", 2245 => "0001010000110100", 2246 => "1101100100001011", 2247 => "0000110000011111", 2248 => "1110010100110100", 2249 => "0100101110111010", 2250 => "1101111110011011", 2251 => "1101101011100011", 2252 => "0010000001010011", 2253 => "1011000000011111", 2254 => "1011010001001001", 2255 => "0100111000100111", 2256 => "0010100000101111", 2257 => "0011101010011101", 2258 => "0010110010111010", 2259 => "1011111110111011", 2260 => "1011010100011010", 2261 => "0101110010101111", 2262 => "0111011111100101", 2263 => "0000010101101110", 2264 => "1011111110001100", 2265 => "1111011101101100", 2266 => "1101011101111000", 2267 => "0010011110000010", 2268 => "0100100000010001", 2269 => "0110010111000011", 2270 => "1110111101011000", 2271 => "0001100110000010", 2272 => "0010001111010011", 2273 => "0111001110110011", 2274 => "1111100100000010", 2275 => "0110101110000011", 2276 => "1000100011100000", 2277 => "1110100101101001", 2278 => "0010000110100110", 2279 => "1101001101001110", 2280 => "0000011011010110", 2281 => "0111101001101110", 2282 => "1101110101111101", 2283 => "0110000010101110", 2284 => "0001000011101111", 2285 => "1100100100110111", 2286 => "1100110111101110", 2287 => "0011010000111000", 2288 => "1010111011011110", 2289 => "1110000100110111", 2290 => "1101110011010010", 2291 => "0111001011111000", 2292 => "1111000100010011", 2293 => "1110010110101110", 2294 => "1010110100000001", 2295 => "0100101110110000", 2296 => "0111110100110000", 2297 => "0011011011110000", 2298 => "0110011001010111", 2299 => "0111001001010111", 2300 => "1110100111111111", 2301 => "0101110101010111", 2302 => "0101011111011010", 2303 => "0010000111001000", 2304 => "1011000001001110", 2305 => "0011110111110000", 2306 => "1000010101001110", 2307 => "0110000100000111", 2308 => "1010100000000111", 2309 => "0101110100001011", 2310 => "1110100110100101", 2311 => "1011100100001111", 2312 => "1101111001111100", 2313 => "0111110000110100", 2314 => "0001010111010001", 2315 => "1010000000001000", 2316 => "1110111011010010", 2317 => "0010110011111011", 2318 => "1011111100000000", 2319 => "1100010010001011", 2320 => "0011000011111011", 2321 => "1110111010111100", 2322 => "1001101001110011", 2323 => "0011010100001100", 2324 => "1111001100010110", 2325 => "0111110011111010", 2326 => "0101011010110111", 2327 => "1010010001001001", 2328 => "0001011111101010", 2329 => "1110011100111011", 2330 => "0011010101001110", 2331 => "1011011111011110", 2332 => "0011001010000100", 2333 => "1001001000101010", 2334 => "1010010100010111", 2335 => "1100001110010000", 2336 => "1110010010000100", 2337 => "1101110111111100", 2338 => "1011001001000111", 2339 => "1111010001001100", 2340 => "1110111100001011", 2341 => "1111111010010100", 2342 => "1010011000011101", 2343 => "0001001100110000", 2344 => "1011010011110110", 2345 => "0110110101110100", 2346 => "0111000001001010", 2347 => "1011001100101101", 2348 => "0011010011100110", 2349 => "0001101100001011", 2350 => "1100101101010001", 2351 => "0011011110101001", 2352 => "1101101010101101", 2353 => "1011100010011110", 2354 => "1110110010110101", 2355 => "0001110000000100", 2356 => "1000001101110010", 2357 => "1010100110100100", 2358 => "1001111100011101", 2359 => "1000010001100111", 2360 => "0111010111000000", 2361 => "0001000001111100", 2362 => "0111110100011110", 2363 => "0100101101111010", 2364 => "0000111111011110", 2365 => "0010001111001000", 2366 => "1100011110111110", 2367 => "0000001001101111", 2368 => "0010001001000001", 2369 => "0111000001111001", 2370 => "0110000101011011", 2371 => "1000101000010110", 2372 => "1100001001100001", 2373 => "0010110000011111", 2374 => "0110111111000101", 2375 => "1100111101001010", 2376 => "0000010010111010", 2377 => "1101000101000101", 2378 => "0110101111010000", 2379 => "0101111110011110", 2380 => "1000011011000010", 2381 => "0101010110000001", 2382 => "0111110001101010", 2383 => "0100111000100011", 2384 => "0011101011011000", 2385 => "0110000011010010", 2386 => "1111010101011111", 2387 => "1000000111011011", 2388 => "0001101100010001", 2389 => "1111111011101010", 2390 => "1010111010111011", 2391 => "1000111110100110", 2392 => "0111100111101110", 2393 => "0100101001001100", 2394 => "0011000100001101", 2395 => "1101100011000011", 2396 => "0100101011100110", 2397 => "0010000110101110", 2398 => "1100010101110001", 2399 => "1001001111110100", 2400 => "1000110001010110", 2401 => "1110001101110010", 2402 => "1110011010010011", 2403 => "0100001010111001", 2404 => "1111011001100010", 2405 => "1000111100011010", 2406 => "0111110100111101", 2407 => "0011010010000110", 2408 => "0011001110001101", 2409 => "1011111100010001", 2410 => "0000001100101010", 2411 => "1100010110111110", 2412 => "1110010110001111", 2413 => "0010100101000111", 2414 => "1110010000110101", 2415 => "1100000111010110", 2416 => "0101101001011101", 2417 => "1001111010100101", 2418 => "1001000110101110", 2419 => "1010100100010100", 2420 => "0101000011111001", 2421 => "0110101001010001", 2422 => "1000100001010001", 2423 => "0000111000101110", 2424 => "1100001010010101", 2425 => "1101110010110000", 2426 => "0001001111000101", 2427 => "1000000001011110", 2428 => "1100011000100100", 2429 => "1100101111110101", 2430 => "1100011011110110", 2431 => "1110110101010100", 2432 => "1101100001110110", 2433 => "0011011010110110", 2434 => "1100110100110110", 2435 => "0000001001111001", 2436 => "0010011011000000", 2437 => "1001010011111001", 2438 => "0001001101100110", 2439 => "1110010011001010", 2440 => "0100001111011111", 2441 => "0011011000100110", 2442 => "1110110011011110", 2443 => "1101001000100001", 2444 => "0001000000000011", 2445 => "0100011100111000", 2446 => "1011010010000101", 2447 => "1000010111101000", 2448 => "0111000101000000", 2449 => "1010011111110010", 2450 => "0101111101000001", 2451 => "0110011100000100", 2452 => "0000111001111011", 2453 => "0010111000110100", 2454 => "1010100010101000", 2455 => "0100001110101111", 2456 => "1110111010110111", 2457 => "1000100110011111", 2458 => "0011110101010110", 2459 => "0111100010100001", 2460 => "0101111010001110", 2461 => "0001000100111110", 2462 => "1100010000110111", 2463 => "0000000010101100", 2464 => "1101101100101011", 2465 => "0000111110001110", 2466 => "0111101100111101", 2467 => "1100010110001000", 2468 => "0111001110011100", 2469 => "0111100111010101", 2470 => "1100000110001111", 2471 => "0101100111101010", 2472 => "1111101111111011", 2473 => "1111001101100011", 2474 => "0110000010111101", 2475 => "0110100000110100", 2476 => "0011011110100100", 2477 => "0100110010101010", 2478 => "1011110001110110", 2479 => "1000101101101011", 2480 => "0111011000001111", 2481 => "1010111110111110", 2482 => "0110011010011010", 2483 => "1000111101010001", 2484 => "1010010001001101", 2485 => "1111110001001110", 2486 => "0111101111001000", 2487 => "0101111111011100", 2488 => "0011001010101100", 2489 => "1100000110000100", 2490 => "0110010111100111", 2491 => "1000110000011110", 2492 => "0111001101010110", 2493 => "1111101011010000", 2494 => "1001111111001110", 2495 => "0111111101010110", 2496 => "0111000001110100", 2497 => "1101111000110001", 2498 => "0000000011110110", 2499 => "0101100011001000", 2500 => "1001010101110011", 2501 => "0101011010111101", 2502 => "1000011101010111", 2503 => "0110110010010010", 2504 => "1001111010011101", 2505 => "0010111011010000", 2506 => "0011000001001111", 2507 => "1111011000001001", 2508 => "0001001010001010", 2509 => "0000110001000110", 2510 => "1011011001111011", 2511 => "1001111101010101", 2512 => "0000100010110111", 2513 => "0111000110010000", 2514 => "0101001101111001", 2515 => "1000111101011111", 2516 => "1101110100110100", 2517 => "0100100000101001", 2518 => "1001111101101110", 2519 => "1010101101011010", 2520 => "1110001011100101", 2521 => "1001010010110011", 2522 => "1010010001010111", 2523 => "0011100001101110", 2524 => "1011000000111011", 2525 => "1101101010111101", 2526 => "0110001000110001", 2527 => "0101100000110001", 2528 => "0010011010000101", 2529 => "0110110000110000", 2530 => "1110001101111000", 2531 => "1100000011000111", 2532 => "1000001000011100", 2533 => "0110101000010101", 2534 => "1111000001100101", 2535 => "1110100001011110", 2536 => "0100001000111001", 2537 => "1000011100000100", 2538 => "0101111000010111", 2539 => "1000110000000000", 2540 => "1011101011110001", 2541 => "0011010000001001", 2542 => "0101101101010000", 2543 => "1100000101101001", 2544 => "0000010101100000", 2545 => "1100100010010111", 2546 => "1010100011100010", 2547 => "1001010110111010", 2548 => "1111000011010100", 2549 => "0000000110011100", 2550 => "0111110111000111", 2551 => "1100111100011001", 2552 => "1000111000000100", 2553 => "0001111001010110", 2554 => "1011001110010001", 2555 => "1110100000001100", 2556 => "1010100101001001", 2557 => "1010000110100110", 2558 => "0101011111010010", 2559 => "1111111010010011", 2560 => "0101011000101001", 2561 => "1111101111101111", 2562 => "1010110000100110", 2563 => "1001000111110100", 2564 => "0011011110111001", 2565 => "1001111001011000", 2566 => "1101010111001111", 2567 => "0101011100011001", 2568 => "1100000101000001", 2569 => "1010110001011000", 2570 => "1001011010011000", 2571 => "0000110101011000", 2572 => "0001111100011111", 2573 => "0111010111110011", 2574 => "0101110010000001", 2575 => "1100010101001110", 2576 => "0100000010011101", 2577 => "0110111010111001", 2578 => "1111100100110111", 2579 => "1010011011010100", 2580 => "1100000010110000", 2581 => "1100010010010110", 2582 => "1011100010000011", 2583 => "0100000010111011", 2584 => "1110110111000100", 2585 => "0010001010100101", 2586 => "1100100101000101", 2587 => "1011011111110101", 2588 => "0010000010010011", 2589 => "1111101000101111", 2590 => "1111111110101001", 2591 => "0010110110101110", 2592 => "1010110101010010", 2593 => "0001001100001101", 2594 => "1000011010001110", 2595 => "1000110001100111", 2596 => "0001111100110100", 2597 => "0010001010010000", 2598 => "1001110000011111", 2599 => "1000001101111011", 2600 => "0011011011011100", 2601 => "1010011010000110", 2602 => "0110111110000011", 2603 => "0100010011001101", 2604 => "1011100100001000", 2605 => "1111011101100111", 2606 => "1010101000111010", 2607 => "1010100101101001", 2608 => "1100011111011011", 2609 => "1110000101110100", 2610 => "0000111001010000", 2611 => "1001100100100101", 2612 => "1111001110010110", 2613 => "0011111010001010", 2614 => "1000010100101110", 2615 => "0100111001001110", 2616 => "1100100000001111", 2617 => "1100111000001110", 2618 => "1111011000111010", 2619 => "1010000011000110", 2620 => "1011100100100100", 2621 => "0101101000011100", 2622 => "1000101100100100", 2623 => "1001000111110000", 2624 => "1011111100000111", 2625 => "1011110011111110", 2626 => "1111011101110111", 2627 => "1001111010110100", 2628 => "1100000111011010", 2629 => "1111011000011010", 2630 => "0011101111101001", 2631 => "1010000010101100", 2632 => "0110010100001010", 2633 => "0100100111011111", 2634 => "0011100001011101", 2635 => "1100100101000101", 2636 => "1010110001110000", 2637 => "1111011011000011", 2638 => "1011000110111000", 2639 => "1100000000010101", 2640 => "0000001100001000", 2641 => "1100111100010111", 2642 => "0000101000010001", 2643 => "0111001100111000", 2644 => "0010110011111001", 2645 => "0101001110010111", 2646 => "0000101010110001", 2647 => "0110101011011010", 2648 => "1001110101010110", 2649 => "1011111110111001", 2650 => "1101111011100001", 2651 => "1101001010111000", 2652 => "0100110001011110", 2653 => "0010011000001111", 2654 => "1010100100001111", 2655 => "1111000100101000", 2656 => "1010101101100110", 2657 => "0000001111011010", 2658 => "0110111111100010", 2659 => "0111001100000001", 2660 => "1101101101100001", 2661 => "1000100010111111", 2662 => "1000011000000001", 2663 => "0100100010010010", 2664 => "1100001111101000", 2665 => "0000010110111101", 2666 => "0110001011111100", 2667 => "0011000010111000", 2668 => "0111111011000010", 2669 => "0100000000111010", 2670 => "1001011101110111", 2671 => "1011010010100000", 2672 => "1011010111000110", 2673 => "0011100000000110", 2674 => "1111011100000101", 2675 => "0010011001010110", 2676 => "0011010111001111", 2677 => "0001001110100101", 2678 => "0010111111110111", 2679 => "0111000101010101", 2680 => "0110111101011001", 2681 => "0101001110100001", 2682 => "0010010100110100", 2683 => "0110100011001111", 2684 => "1111001000000101", 2685 => "0001001111101100", 2686 => "0001100011100110", 2687 => "1110111100101111", 2688 => "1111011101110100", 2689 => "0101100000000110", 2690 => "0011101101000000", 2691 => "0110000100110111", 2692 => "0111011010111010", 2693 => "0101100001100011", 2694 => "0010010000111111", 2695 => "1011111011011010", 2696 => "0110111000101000", 2697 => "0000010111001001", 2698 => "0000001101100001", 2699 => "0110011001010011", 2700 => "0001110000110011", 2701 => "1011000111100111", 2702 => "0010001101101111", 2703 => "0100010001100110", 2704 => "1110101111100111", 2705 => "0010110000100110", 2706 => "0100101011101101", 2707 => "1011101101101101", 2708 => "1000011100010010", 2709 => "1111100110101100", 2710 => "0100110000011001", 2711 => "1001000101111001", 2712 => "1100001000010010", 2713 => "1010100101111100", 2714 => "0001111110111111", 2715 => "0000001101010100", 2716 => "0100001111101011", 2717 => "0001101101111101", 2718 => "0000011001110110", 2719 => "1010100000110011", 2720 => "0111101011010100", 2721 => "0110101011000110", 2722 => "0100110100011110", 2723 => "0001010000011011", 2724 => "0000101110000001", 2725 => "1111111010011001", 2726 => "0111010001011111", 2727 => "0110000110101111", 2728 => "1001000001011101", 2729 => "1001011000011000", 2730 => "0111101101100110", 2731 => "0110101001110100", 2732 => "1001100111101010", 2733 => "1000111111100100", 2734 => "1001000100000110", 2735 => "0101001010100000", 2736 => "0001011011011100", 2737 => "0101100000110001", 2738 => "0000010000001010", 2739 => "0111111010101110", 2740 => "1100001111111000", 2741 => "0100110110011011", 2742 => "1001101100010001", 2743 => "0110000101010101", 2744 => "1101100110110110", 2745 => "0011000011001110", 2746 => "0000100011000100", 2747 => "0000001100011001", 2748 => "0010011000111100", 2749 => "1110110110000111", 2750 => "1100110001100111", 2751 => "0011001100110011", 2752 => "0111111001001001", 2753 => "1100111101111111", 2754 => "1001111111010010", 2755 => "1111110110111001", 2756 => "0110010100101010", 2757 => "1001011010011001", 2758 => "1111001100000001", 2759 => "1101111000111101", 2760 => "1000011011110000", 2761 => "0111101101010000", 2762 => "0011001101110011", 2763 => "0110001010110000", 2764 => "1011111111001111", 2765 => "1110111110110111", 2766 => "1001111001101000", 2767 => "0001010100110011", 2768 => "0101100010101000", 2769 => "0101101010101100", 2770 => "0110011000110100", 2771 => "0010111001110101", 2772 => "0001110110111111", 2773 => "0110010000100001", 2774 => "1010001001000111", 2775 => "0001000011101011", 2776 => "1010011100100101", 2777 => "0111100010111000", 2778 => "1000111000110100", 2779 => "0000001101010000", 2780 => "0100011000111011", 2781 => "0011011100011111", 2782 => "1000110010101011", 2783 => "0101101110111110", 2784 => "1010111110100011", 2785 => "1110101101101100", 2786 => "1011101010011110", 2787 => "1001011000111011", 2788 => "1010101111100100", 2789 => "1011010101111111", 2790 => "1001101100111011", 2791 => "1100000100101100", 2792 => "0100101100000110", 2793 => "1100111100110111", 2794 => "1011001111011101", 2795 => "0000110100011001", 2796 => "0011100111101001", 2797 => "1001110110110101", 2798 => "1111001101110000", 2799 => "0001011010100110", 2800 => "0000011110001110", 2801 => "1111101100111001", 2802 => "1000010001111010", 2803 => "1101001100111011", 2804 => "1100000110110010", 2805 => "0010001011001101", 2806 => "1011100110101111", 2807 => "0100000100001100", 2808 => "1011111100100101", 2809 => "0111100100111101", 2810 => "0101001001100011", 2811 => "1100101001110111", 2812 => "0000001111010100", 2813 => "0111001011010001", 2814 => "0001100000010100", 2815 => "1111011010101001", 2816 => "1101101000011100", 2817 => "1011100110111101", 2818 => "1111101001010101", 2819 => "0000111110111011", 2820 => "1001111111010101", 2821 => "0001110000000001", 2822 => "1011101001011010", 2823 => "0001111101000101", 2824 => "1001001111000010", 2825 => "1000000111100110", 2826 => "0000100101010100", 2827 => "1101010101010000", 2828 => "1011000100011001", 2829 => "0101011000001010", 2830 => "0000010000100001", 2831 => "1101100111110010", 2832 => "0101010001000001", 2833 => "1001010101100100", 2834 => "1100011000000111", 2835 => "0110000101100010", 2836 => "0000100001110010", 2837 => "0110011011010111", 2838 => "0011000110101111", 2839 => "0001001000110111", 2840 => "1100010010101100", 2841 => "0010001100011100", 2842 => "1010000101001111", 2843 => "1010111111101001", 2844 => "1011110101010100", 2845 => "0000110010001100", 2846 => "0010011101110101", 2847 => "1011001111101010", 2848 => "0101101100111011", 2849 => "1100000011010001", 2850 => "1001110000111111", 2851 => "1101100111001100", 2852 => "0110000010100010", 2853 => "1110000010110000", 2854 => "0001110001011000", 2855 => "0010000011110100", 2856 => "1101111110010110", 2857 => "0101011001111111", 2858 => "0000010001100000", 2859 => "1111011111110100", 2860 => "1000001101001010", 2861 => "0010001100000101", 2862 => "1001110111101111", 2863 => "1110000100111011", 2864 => "1100111011101001", 2865 => "0101101110000011", 2866 => "1101100010000101", 2867 => "0011001000101111", 2868 => "1110001011011001", 2869 => "0000101010001110", 2870 => "0000000010010110", 2871 => "1110111101010110", 2872 => "0111000010001011", 2873 => "1111011101000010", 2874 => "1101001010101101", 2875 => "0011110111000011", 2876 => "0000101101000001", 2877 => "0100000000101100", 2878 => "1010010010100000", 2879 => "1001100001011101", 2880 => "1101000101000011", 2881 => "0000100111010110", 2882 => "0001011111110000", 2883 => "1111110000001111", 2884 => "0111011100101001", 2885 => "0100110001000100", 2886 => "0111100100111100", 2887 => "1001010001111110", 2888 => "0010011010011111", 2889 => "0010111010100000", 2890 => "0011101010001111", 2891 => "1000011010110101", 2892 => "1000110101111011", 2893 => "0111001010100110", 2894 => "1101011001010010", 2895 => "1011101111010000", 2896 => "0111110010000001", 2897 => "1101111101011100", 2898 => "0000111101111110", 2899 => "0011001011101101", 2900 => "0101110010001100", 2901 => "0110100101111010", 2902 => "0101001100011001", 2903 => "0010011001001110", 2904 => "1110011101111011", 2905 => "1001110001010000", 2906 => "0001101010000001", 2907 => "1011100000000100", 2908 => "1100011111010110", 2909 => "1011100010110000", 2910 => "1110100101110101", 2911 => "0100111110001110", 2912 => "0000100000110011", 2913 => "0010001001111011", 2914 => "0100101100110001", 2915 => "0100010100110011", 2916 => "1010110010000101", 2917 => "0100111110111000", 2918 => "1111100100100111", 2919 => "0010010100000110", 2920 => "1010110111000111", 2921 => "1011100101001101", 2922 => "1100001101010101", 2923 => "1010100101001011", 2924 => "0100010111000101", 2925 => "1000101110000100", 2926 => "1010011100011100", 2927 => "1100110100001101", 2928 => "1111011010110010", 2929 => "1001011100010010", 2930 => "0101000001101000", 2931 => "1000011111011000", 2932 => "0100110011000010", 2933 => "1011011110011100", 2934 => "1110110000101111", 2935 => "0110100000001011", 2936 => "0000100000011001", 2937 => "1110000111001001", 2938 => "0001110010001000", 2939 => "1000110001100011", 2940 => "0010101111111101", 2941 => "1101011111110111", 2942 => "0011001010010111", 2943 => "0001011000010101", 2944 => "1000010100001001", 2945 => "0110110001010011", 2946 => "1000101111000010", 2947 => "0001111111100110", 2948 => "1100011010010100", 2949 => "0110101101000110", 2950 => "1001001010011100", 2951 => "0000000001010010", 2952 => "1001010101111011", 2953 => "1100111000001011", 2954 => "1001000110010111", 2955 => "1000011001011101", 2956 => "0011001000100000", 2957 => "1101110101100111", 2958 => "0110011111011100", 2959 => "0001111110100101", 2960 => "1010001101100011", 2961 => "0010000000101010", 2962 => "0010010100000110", 2963 => "0100000111000010", 2964 => "1110001110101001", 2965 => "0110011101001011", 2966 => "0110111000000111", 2967 => "0001011110000110", 2968 => "1001001010110000", 2969 => "1110101100000111", 2970 => "1010000111101001", 2971 => "0101111000100111", 2972 => "0111110110000010", 2973 => "1001100101010010", 2974 => "0001110000011110", 2975 => "1010100101001011", 2976 => "0010011111010001", 2977 => "1101010100001000", 2978 => "1111101101000010", 2979 => "0011001101110011", 2980 => "1100000111010101", 2981 => "0011011100101111", 2982 => "0111111110101101", 2983 => "0110010110101010", 2984 => "0010001110111011", 2985 => "1011101101100010", 2986 => "0110111010110011", 2987 => "1000111000100011", 2988 => "0011011100000101", 2989 => "0001011010110101", 2990 => "1000011101001000", 2991 => "0101001000001111", 2992 => "1110101111111110", 2993 => "1100011101000101", 2994 => "0101111000111000", 2995 => "1011100111101111", 2996 => "0010011111001111", 2997 => "1001101101000010", 2998 => "1010111111010111", 2999 => "0101000111111010", 3000 => "0011110110110100", 3001 => "1110111100001010", 3002 => "0101000000010110", 3003 => "0010101011000000", 3004 => "0010000000011100", 3005 => "1110111000010101", 3006 => "1000111110110101", 3007 => "0101011011110001", 3008 => "1111011100001111", 3009 => "1001111000110110", 3010 => "0111011100110001", 3011 => "0101110100111110", 3012 => "0001000001001000", 3013 => "0001100011010100", 3014 => "0001110111111010", 3015 => "1101001011100000", 3016 => "0100000010110101", 3017 => "1000101011100010", 3018 => "0000101111111110", 3019 => "1101110101010000", 3020 => "0100011101111110", 3021 => "1100111010011010", 3022 => "1111010111010101", 3023 => "1100111010111110", 3024 => "0111011110111101", 3025 => "0100001010000001", 3026 => "1000111010101101", 3027 => "0110000001011101", 3028 => "1111110110011001", 3029 => "0010100001001000", 3030 => "1010011010100100", 3031 => "0101110011110111", 3032 => "1100101000111000", 3033 => "0010001010011011", 3034 => "0110110000101110", 3035 => "1001110001111000", 3036 => "0100100010111111", 3037 => "1101101010001111", 3038 => "0100101000101110", 3039 => "1111101101100000", 3040 => "1000000111111100", 3041 => "1101110010111001", 3042 => "1111101001110101", 3043 => "0000000110010001", 3044 => "0011000110110100", 3045 => "1001000001101111", 3046 => "1101101110010111", 3047 => "0111110100100001", 3048 => "1011011000110101", 3049 => "0110101000101010", 3050 => "0000000100000101", 3051 => "0010111011011110", 3052 => "0111001111110011", 3053 => "1110010001101101", 3054 => "0001110011101110", 3055 => "0011001001000100", 3056 => "0000001000010010", 3057 => "1100110010001110", 3058 => "0010000000010111", 3059 => "1111100001000001", 3060 => "0100101000100011", 3061 => "1101110111000000", 3062 => "1011000001100000", 3063 => "1000011011111001", 3064 => "0010110111101010", 3065 => "1001110101011110", 3066 => "1000110011000001", 3067 => "1000110110110000", 3068 => "1001000001111011", 3069 => "1110010100101001", 3070 => "0000001010000011", 3071 => "1111101101011010", 3072 => "1100000001000001", 3073 => "1100110011101100", 3074 => "1110111011001110", 3075 => "0010000101011001", 3076 => "1000000000000000", 3077 => "1100110100000010", 3078 => "0100111000110010", 3079 => "1100011111000111", 3080 => "1100011000000011", 3081 => "0000100001011000", 3082 => "0001010010000011", 3083 => "1010110000011101", 3084 => "0111110010011011", 3085 => "1100011101110000", 3086 => "0001000100000111", 3087 => "1110101101110010", 3088 => "1111000001100010", 3089 => "1100010101000000", 3090 => "1111010010100101", 3091 => "1000001101000101", 3092 => "0100011011100010", 3093 => "1110101011110010", 3094 => "1100101100110000", 3095 => "1011100100010101", 3096 => "1110011100001111", 3097 => "1111010001101100", 3098 => "0110111100101001", 3099 => "1100000000111111", 3100 => "1000100101110111", 3101 => "0011001100101101", 3102 => "1011010111110110", 3103 => "0101100110010001", 3104 => "1001100111100100", 3105 => "0011100001010110", 3106 => "0001010001100100", 3107 => "0101001010111101", 3108 => "0011111100110010", 3109 => "1010100101101011", 3110 => "0001100110010001", 3111 => "1100110101111011", 3112 => "0100011100110111", 3113 => "0100110000000101", 3114 => "1000111000101001", 3115 => "0010101100010101", 3116 => "1011111010011110", 3117 => "0100100000011000", 3118 => "1010001100011101", 3119 => "1111100010010110", 3120 => "1010010000110101", 3121 => "0001110111000110", 3122 => "1010101001110010", 3123 => "0010001010101111", 3124 => "0000001011000100", 3125 => "0110101101101000", 3126 => "1110010011000111", 3127 => "0100101100011111", 3128 => "1111101111001100", 3129 => "1110011000111110", 3130 => "0101100100001100", 3131 => "1110010100101000", 3132 => "0011011010110000", 3133 => "0010100011100001", 3134 => "1110001010001000", 3135 => "0010100010110101", 3136 => "0101001110101100", 3137 => "0011110011110110", 3138 => "1111100011000010", 3139 => "1010010010100001", 3140 => "0100100001011111", 3141 => "1000110001111111", 3142 => "0001000011001010", 3143 => "1011110000110001", 3144 => "1111001110010001", 3145 => "1111011100110001", 3146 => "1001110110110111", 3147 => "0101000011011110", 3148 => "0011011011001111", 3149 => "0011000000010001", 3150 => "1001000101001001", 3151 => "1001000010111010", 3152 => "0101100010001110", 3153 => "0100110110011111", 3154 => "0101100110010000", 3155 => "1010110100000110", 3156 => "0001011110111011", 3157 => "1001011010010101", 3158 => "0011000011111100", 3159 => "1001011011101011", 3160 => "1110010011100111", 3161 => "1101000100100010", 3162 => "1111100101100001", 3163 => "0111100100010100", 3164 => "1100000100001110", 3165 => "1000110110100010", 3166 => "1111110001000101", 3167 => "1001001110010000", 3168 => "0010001100100001", 3169 => "0101010101011111", 3170 => "1000101000001011", 3171 => "0000000011101000", 3172 => "1011101011101011", 3173 => "1010111101110001", 3174 => "0111000011110101", 3175 => "0000110001101011", 3176 => "0000101100001010", 3177 => "1011100101000100", 3178 => "0011101010001100", 3179 => "0011001011000101", 3180 => "1001111010101001", 3181 => "1101011111101011", 3182 => "1110111000101010", 3183 => "1011000000001010", 3184 => "0110110111001101", 3185 => "1100001000010001", 3186 => "0010100001000000", 3187 => "0111110010100010", 3188 => "0111100111010110", 3189 => "1010111000010100", 3190 => "0011110110100110", 3191 => "1110110110100101", 3192 => "1010111001110101", 3193 => "0100110011101100", 3194 => "1000010100011101", 3195 => "1111100101000100", 3196 => "1000110110110010", 3197 => "1011011101111000", 3198 => "1010110110010111", 3199 => "0111001101000101", 3200 => "0110000110101110", 3201 => "1111010001010111", 3202 => "0100001100011111", 3203 => "1001001110011111", 3204 => "1011110011001101", 3205 => "1110110000001011", 3206 => "0001011010111000", 3207 => "0010101011010010", 3208 => "0100010101011111", 3209 => "0111011111001110", 3210 => "0100111111111110", 3211 => "0111010100110110", 3212 => "1011010111010000", 3213 => "1000000011110101", 3214 => "0110000110110010", 3215 => "0101100010011010", 3216 => "0111000100100010", 3217 => "0001111100011010", 3218 => "0101010011101001", 3219 => "1011110010011001", 3220 => "0100010010100100", 3221 => "1110100010000110", 3222 => "0100000011111111", 3223 => "0111001001111001", 3224 => "1110100111010011", 3225 => "1110010010001101", 3226 => "0111100000110110", 3227 => "1010100010011010", 3228 => "1101001010001000", 3229 => "1111110010101111", 3230 => "1000110111101111", 3231 => "1110001110100100", 3232 => "1101101010100111", 3233 => "0111111000110101", 3234 => "0110011011010011", 3235 => "1100111000001110", 3236 => "0110111000110010", 3237 => "1000100111100110", 3238 => "1111000111010100", 3239 => "0010100101111001", 3240 => "0101100100101110", 3241 => "1101110100000100", 3242 => "0111110100000001", 3243 => "1011101100010010", 3244 => "1100010001000010", 3245 => "0010001011000110", 3246 => "0110000000110101", 3247 => "1001101001011000", 3248 => "1010001001110011", 3249 => "0010001011010011", 3250 => "0110100011010101", 3251 => "0110101010010010", 3252 => "1101000001101001", 3253 => "0111101011000011", 3254 => "1111101010101101", 3255 => "1100100110011111", 3256 => "0111011101000000", 3257 => "0001110000110101", 3258 => "0011001100111000", 3259 => "0010011010000001", 3260 => "0111010100110000", 3261 => "0110010101101101", 3262 => "1101010100101001", 3263 => "0001011000100010", 3264 => "0111000101101000", 3265 => "0101111101011010", 3266 => "1001010101101110", 3267 => "1011101111001111", 3268 => "1011010001010011", 3269 => "1011111101000100", 3270 => "1001000111110101", 3271 => "0100000001010100", 3272 => "0110001001111100", 3273 => "0010100010000100", 3274 => "0110010000011110", 3275 => "1111101101100100", 3276 => "1010000101100100", 3277 => "0011111101001000", 3278 => "0111100010000100", 3279 => "1001011001010010", 3280 => "1010000010001111", 3281 => "0110010000010100", 3282 => "0111111001100011", 3283 => "0010011110000000", 3284 => "1010011100001010", 3285 => "0010101111111010", 3286 => "0111001100100011", 3287 => "0111110100100011", 3288 => "0101010000000001", 3289 => "0001110110110000", 3290 => "0011110001011111", 3291 => "1100000111100101", 3292 => "1000000011011000", 3293 => "1010001111101101", 3294 => "1101110010101110", 3295 => "0010001100101111", 3296 => "0000110011010101", 3297 => "1000001001000100", 3298 => "0100011111100000", 3299 => "0010100101000011", 3300 => "0111010011110010", 3301 => "0111001010100011", 3302 => "0011001000010000", 3303 => "1001001101011001", 3304 => "0110001000111001", 3305 => "0010100111111111", 3306 => "1010110101111111", 3307 => "0111000101110001", 3308 => "1111011100110001", 3309 => "0000000111010100", 3310 => "1110010110001001", 3311 => "1001000001000110", 3312 => "0110111100101101", 3313 => "1110011010100111", 3314 => "0110000100001111", 3315 => "0000001001010010", 3316 => "1011010111011011", 3317 => "1001110111001011", 3318 => "0101001110101111", 3319 => "0010110011010111", 3320 => "0010001110110011", 3321 => "0001011100011111", 3322 => "1001110011010100", 3323 => "1101101011001001", 3324 => "1111001011000100", 3325 => "1001010100001110", 3326 => "0111000111100010", 3327 => "0110011101100000", 3328 => "1110000011110011", 3329 => "1101010110001110", 3330 => "1101111010010111", 3331 => "0101100101111011", 3332 => "1100101001111001", 3333 => "0101110100000111", 3334 => "1010111101001010", 3335 => "1100010000001001", 3336 => "1011011111011010", 3337 => "1000111000010000", 3338 => "0100000100100010", 3339 => "1101001101100111", 3340 => "0101010010010110", 3341 => "0000011101111001", 3342 => "0011000000100000", 3343 => "1001011001101001", 3344 => "0011101111001010", 3345 => "0100011111110011", 3346 => "1111010101001100", 3347 => "1100010010111011", 3348 => "0011111011001111", 3349 => "0000111111000100", 3350 => "0100100100111000", 3351 => "0011100000101100", 3352 => "1101110111111000", 3353 => "0110110010111100", 3354 => "1001100010111101", 3355 => "1010000010000001", 3356 => "0100011100101100", 3357 => "1011100000111011", 3358 => "0101011100100010", 3359 => "0111010010011000", 3360 => "1001111111101111", 3361 => "1001001000011111", 3362 => "0000111001101011", 3363 => "0110010000100001", 3364 => "0001011101000011", 3365 => "0111111101110100", 3366 => "1101000010100110", 3367 => "0100101000110110", 3368 => "0100001011000111", 3369 => "1101000010111100", 3370 => "1010011011000010", 3371 => "1101100011100110", 3372 => "0100101100101000", 3373 => "0000100011010111", 3374 => "1101110010010000", 3375 => "0110111011010010", 3376 => "1110101010101010", 3377 => "1111000111010000", 3378 => "0110000100001101", 3379 => "1111100111011011", 3380 => "1011110010111001", 3381 => "0000000111011110", 3382 => "0100110001001110", 3383 => "1010100000001100", 3384 => "0010001111111000", 3385 => "0100110110101110", 3386 => "0011111111010100", 3387 => "0011000101101001", 3388 => "1011001000000000", 3389 => "0011000000010111", 3390 => "1100101110000111", 3391 => "1001100100011100", 3392 => "0110010110010101", 3393 => "0010110111011001", 3394 => "1000100000011011", 3395 => "1100011010010101", 3396 => "1011000100101000", 3397 => "0011001111101111", 3398 => "1111001011001000", 3399 => "0010111011100010", 3400 => "1100101101110001", 3401 => "1000100101000000", 3402 => "1100100110101000", 3403 => "1101011110110001", 3404 => "1111110001101000", 3405 => "0101011010001101", 3406 => "1100101001000110", 3407 => "0000011010101001", 3408 => "0010101110111110", 3409 => "1010000110110110", 3410 => "1101101110010010", 3411 => "1001100110111001", 3412 => "1110110001100011", 3413 => "0100001111010010", 3414 => "1011010000010100", 3415 => "0011101100010110", 3416 => "0011011001010001", 3417 => "0001110000011110", 3418 => "1110101010110111", 3419 => "0110010000111111", 3420 => "0010111000011110", 3421 => "1101000110011010", 3422 => "0010111110001010", 3423 => "1100100101110101", 3424 => "1010011001011000", 3425 => "1010101110001010", 3426 => "1110001010001011", 3427 => "1111001000010101", 3428 => "1110110111011010", 3429 => "1110110110100010", 3430 => "0101100100010011", 3431 => "1000100111000010", 3432 => "1110110110000110", 3433 => "1101101110000100", 3434 => "0110000101011101", 3435 => "0101001100100110", 3436 => "1010110100001110", 3437 => "1011000000100011", 3438 => "1010000001001000", 3439 => "1001110101010110", 3440 => "1011110000100110", 3441 => "0011011001100001", 3442 => "1100111101110101", 3443 => "1101100011011010", 3444 => "0111010100000100", 3445 => "1001101001100000", 3446 => "1101100101001101", 3447 => "1011001000000000", 3448 => "1100010110101000", 3449 => "1010111010000000", 3450 => "1011011000111011", 3451 => "1001000011111101", 3452 => "0100001111100100", 3453 => "0111100110101110", 3454 => "0010100010110000", 3455 => "1011001001011111", 3456 => "0101111110110011", 3457 => "0111010110100011", 3458 => "1101111011010100", 3459 => "1100101010100010", 3460 => "1010010100110011", 3461 => "0101100010111101", 3462 => "0001100110101001", 3463 => "1001011100011100", 3464 => "0001010001110110", 3465 => "1110111010110000", 3466 => "0001110011101011", 3467 => "0000111010110010", 3468 => "1111001110010011", 3469 => "0000001001110001", 3470 => "0010010110110111", 3471 => "0000011101111100", 3472 => "1011110101000100", 3473 => "0001101001111100", 3474 => "1011101100101100", 3475 => "1011111110000001", 3476 => "1001111011111001", 3477 => "1010001111000110", 3478 => "0000111111111011", 3479 => "1010001010100000", 3480 => "0011100110111110", 3481 => "0001101110101010", 3482 => "0011100110111010", 3483 => "1000110000011101", 3484 => "1100000011101000", 3485 => "0110101111101111", 3486 => "1100000011110011", 3487 => "0100101110011110", 3488 => "1110010110111001", 3489 => "0011111000000011", 3490 => "0110100100011000", 3491 => "1111110100011111", 3492 => "0111100001111111", 3493 => "0001000011001000", 3494 => "0111001111010100", 3495 => "1101100111100101", 3496 => "1100110101000001", 3497 => "0000101100100010", 3498 => "0001000110010010", 3499 => "0101001110010010", 3500 => "1001010010110101", 3501 => "1111100110111101", 3502 => "0010000110100001", 3503 => "0000110000111010", 3504 => "1010110010011001", 3505 => "0110101100001101", 3506 => "0001000011100010", 3507 => "0011110101011011", 3508 => "0110010000000000", 3509 => "0001001010111110", 3510 => "1001111011001100", 3511 => "1101100111000011", 3512 => "0111100010111000", 3513 => "0100011100110000", 3514 => "0110001110101011", 3515 => "1000000001010010", 3516 => "0111101000101111", 3517 => "0001010101100110", 3518 => "0001100111010100", 3519 => "1101000001011010", 3520 => "1001100111010011", 3521 => "0001011101110001", 3522 => "1110100000000100", 3523 => "1011111001001010", 3524 => "0111100110100001", 3525 => "1011000111000001", 3526 => "1000111010100110", 3527 => "1001101010110010", 3528 => "0001010011011011", 3529 => "1111000111011110", 3530 => "0110101010100100", 3531 => "0111101010000110", 3532 => "1101111001100000", 3533 => "1011111010111000", 3534 => "0110101111111100", 3535 => "1111011001111101", 3536 => "0010010001001101", 3537 => "0000011000010010", 3538 => "0011010111001011", 3539 => "0011100101110001", 3540 => "0111111000101011", 3541 => "0110110111111100", 3542 => "1000011000100000", 3543 => "1010010100000011", 3544 => "0111101100101111", 3545 => "1111001101001111", 3546 => "0111000111110110", 3547 => "1011010101110100", 3548 => "1010001010110100", 3549 => "1111101101101011", 3550 => "0011111101011011", 3551 => "1100000000000110", 3552 => "1110101000000110", 3553 => "0010011101001011", 3554 => "1011100111110011", 3555 => "0100010100000010", 3556 => "0111010000101100", 3557 => "0111100001011101", 3558 => "0100011110101100", 3559 => "1000001000000110", 3560 => "0111101101011011", 3561 => "1111111010101000", 3562 => "1101001111100110", 3563 => "1000000011000011", 3564 => "1110101101011010", 3565 => "1001000001000011", 3566 => "1110001001101011", 3567 => "1111000011000101", 3568 => "0010110010001100", 3569 => "0110010110101111", 3570 => "0000000001101000", 3571 => "1101000110011110", 3572 => "1011110110010100", 3573 => "1001100101101000", 3574 => "0100101001001100", 3575 => "1001011010110111", 3576 => "0010000100100101", 3577 => "1010110010011101", 3578 => "1111000100101010", 3579 => "0000011100011101", 3580 => "0010000010001111", 3581 => "1111111111100110", 3582 => "1101101011000100", 3583 => "1101111011101110", 3584 => "1011011000100100", 3585 => "1111010000001111", 3586 => "1101010000010110", 3587 => "1000111010010000", 3588 => "1011110101101010", 3589 => "1000101001110001", 3590 => "0010111011100010", 3591 => "1001111101110101", 3592 => "1110111000100010", 3593 => "1001000100011111", 3594 => "1110010100111100", 3595 => "0011101111001100", 3596 => "0111000111100100", 3597 => "0111111100001010", 3598 => "1110001010110010", 3599 => "0010101111100101", 3600 => "1101100101111110", 3601 => "1111111000100000", 3602 => "0110101101000110", 3603 => "0011010011100100", 3604 => "0000110110000000", 3605 => "1000100011111110", 3606 => "1010101011100011", 3607 => "0000000110011110", 3608 => "1100000000110101", 3609 => "1101111100010001", 3610 => "1011001111101111", 3611 => "0110000001010110", 3612 => "1111010101110101", 3613 => "1011100011100100", 3614 => "0001100010001100", 3615 => "1001001011100001", 3616 => "0001110010000000", 3617 => "1000111010010110", 3618 => "1010001001110001", 3619 => "0001100011110001", 3620 => "0101111110111100", 3621 => "1001011111000110", 3622 => "1100000001001000", 3623 => "0011111101001010", 3624 => "1011011001101000", 3625 => "1111011110000111", 3626 => "1100011011011011", 3627 => "1111000010011011", 3628 => "1001010101110000", 3629 => "0011101110101100", 3630 => "0011001111001001", 3631 => "0110001110100100", 3632 => "1010101111011010", 3633 => "1000011000110011", 3634 => "0110001100111101", 3635 => "0111000010011000", 3636 => "0000111111101001", 3637 => "1100011000010010", 3638 => "0001100000110101", 3639 => "0011000110001011", 3640 => "0011000111010010", 3641 => "0011111110011100", 3642 => "1011101000010101", 3643 => "1101011111000011", 3644 => "0111111001111000", 3645 => "0101000110001000", 3646 => "1000000010101011", 3647 => "1011110110011100", 3648 => "0010010100111000", 3649 => "1100111110001101", 3650 => "0101001110001010", 3651 => "0001011000001001", 3652 => "1100111110101110", 3653 => "0100011111111010", 3654 => "0010001011110101", 3655 => "0010001001100001", 3656 => "1010010111101010", 3657 => "0111000100101011", 3658 => "0101000001001001", 3659 => "1010001111000010", 3660 => "0011101010010111", 3661 => "0001010001011100", 3662 => "0110101111110001", 3663 => "1000011110110011", 3664 => "1110111001010000", 3665 => "1011101000110001", 3666 => "1100001010101011", 3667 => "1010001101000111", 3668 => "0001110011111000", 3669 => "0011111111110100", 3670 => "0111101000000000", 3671 => "0111111101000010", 3672 => "1111000110011110", 3673 => "1010000001011010", 3674 => "1011010000101010", 3675 => "1111101000110111", 3676 => "0010011110000000", 3677 => "0111010100011101", 3678 => "0001010000111101", 3679 => "0110001111011010", 3680 => "1101010100011101", 3681 => "0000000001110011", 3682 => "1000110110011000", 3683 => "1000101010101111", 3684 => "1001001000101100", 3685 => "0010101110111000", 3686 => "1110110010000110", 3687 => "0011010010000111", 3688 => "1011001000100000", 3689 => "1000111101110111", 3690 => "0010100011010000", 3691 => "1010110110001000", 3692 => "0110101110111000", 3693 => "0010110000111100", 3694 => "0111110111010111", 3695 => "0100100001010010", 3696 => "0111100100001101", 3697 => "0011000000100001", 3698 => "0111100101101111", 3699 => "1000001101101000", 3700 => "1010000001111011", 3701 => "0001100110100111", 3702 => "0111111010011110", 3703 => "1001111100000010", 3704 => "1010010010100101", 3705 => "0000110011011001", 3706 => "1111011011101001", 3707 => "1001001110011011", 3708 => "0011010001111110", 3709 => "1110010111111111", 3710 => "0101010011000001", 3711 => "1110100110001011", 3712 => "0101001101001000", 3713 => "0010011100010000", 3714 => "1011000001100001", 3715 => "1111111111011110", 3716 => "1010010001100001", 3717 => "0110001111001000", 3718 => "1010110011111100", 3719 => "1011111011000001", 3720 => "0111111001100110", 3721 => "1101101100010000", 3722 => "1101011101000110", 3723 => "0000110011110101", 3724 => "1001111000000011", 3725 => "1001000100111011", 3726 => "1101000001101111", 3727 => "1000111001001111", 3728 => "0010011110010000", 3729 => "1010110000010000", 3730 => "0101001011111000", 3731 => "1011011111111110", 3732 => "0101110000001011", 3733 => "0011101000101011", 3734 => "0100000101000001", 3735 => "1011010110101001", 3736 => "1111110100101010", 3737 => "0100111011110011", 3738 => "0100101110000011", 3739 => "1000110110100000", 3740 => "0110010001011000", 3741 => "1100111010110111", 3742 => "0111001001101001", 3743 => "0110010001101010", 3744 => "0101111101011000", 3745 => "1111001111110000", 3746 => "1110100010001101", 3747 => "1001011101111010", 3748 => "1000000100010111", 3749 => "1100001110010010", 3750 => "1011100100101001", 3751 => "0101101001111010", 3752 => "0110001111000000", 3753 => "1111110000111100", 3754 => "0100101100011101", 3755 => "1111000101001011", 3756 => "1101100100100111", 3757 => "1001110110111100", 3758 => "1010011100010010", 3759 => "1101010011110101", 3760 => "1101000011011110", 3761 => "0010011111011101", 3762 => "1100011101101110", 3763 => "1010000011100001", 3764 => "1010110001001001", 3765 => "1101100110110101", 3766 => "1011111110100110", 3767 => "0110110010000111", 3768 => "0100101101101001", 3769 => "0111111110001000", 3770 => "0001010110110000", 3771 => "1011000000001100", 3772 => "1011110001111001", 3773 => "0000000010000000", 3774 => "1101011010100100", 3775 => "1011111111010101", 3776 => "0100001111101101", 3777 => "1001010111110110", 3778 => "1010111100000111", 3779 => "1110110011000111", 3780 => "1101111011111010", 3781 => "0011011101010010", 3782 => "1101011111111100", 3783 => "0001110011000101", 3784 => "0001001011100011", 3785 => "1010101001110111", 3786 => "0101000000001001", 3787 => "0100101101101111", 3788 => "1110110111111111", 3789 => "1010011111001011", 3790 => "0101100110100111", 3791 => "0111010001010110", 3792 => "0010100011110110", 3793 => "0001110011010000", 3794 => "1011111000101001", 3795 => "0000101010111010", 3796 => "1000111111100011", 3797 => "0001010101110010", 3798 => "0010001001110010", 3799 => "0110000000100001", 3800 => "1000000010011101", 3801 => "1001010011011101", 3802 => "1000011001111000", 3803 => "0001001011100110", 3804 => "1111100111000001", 3805 => "1011100000010000", 3806 => "1111111100111000", 3807 => "0000100011101011", 3808 => "1011010100111010", 3809 => "1011111010010110", 3810 => "1101001010010011", 3811 => "1011100101110111", 3812 => "0110100101110010", 3813 => "0110000101110101", 3814 => "0011001101111100", 3815 => "1110001110100111", 3816 => "1101110000110011", 3817 => "1010111000010110", 3818 => "1110001001011110", 3819 => "0010111111000010", 3820 => "0000110100101010", 3821 => "0001111110010000", 3822 => "1010001101100001", 3823 => "1011001111001110", 3824 => "1001110110000011", 3825 => "1110000111101101", 3826 => "0100011101101010", 3827 => "0101000110010101", 3828 => "0101111111001101", 3829 => "0011010100001100", 3830 => "0011000111001111", 3831 => "1011011100101111", 3832 => "1010110101110110", 3833 => "1010001010001110", 3834 => "0010001000100000", 3835 => "0111011111110111", 3836 => "1001111110100000", 3837 => "0000011100010000", 3838 => "0010000101110101", 3839 => "0101010011111001", 3840 => "1000101111010001", 3841 => "0000110011101110", 3842 => "0100111101101101", 3843 => "0101000000111010", 3844 => "0011100010001010", 3845 => "0000001100110000", 3846 => "1101111001101101", 3847 => "0011010101100101", 3848 => "0001101001100000", 3849 => "0001000000111100", 3850 => "1111101111011101", 3851 => "1001110011110000", 3852 => "1001101101111011", 3853 => "1111011000100000", 3854 => "1100110100111011", 3855 => "0011111010010101", 3856 => "1100011010010110", 3857 => "1111110110100111", 3858 => "0110111111100011", 3859 => "1000111010010001", 3860 => "1000111111100011", 3861 => "0011001110010111", 3862 => "0111111111100000", 3863 => "1111110100100010", 3864 => "1010001011000001", 3865 => "0110110000100001", 3866 => "0111111111110011", 3867 => "1111111101100100", 3868 => "1110101001100010", 3869 => "1111111101000001", 3870 => "0001001101011111", 3871 => "1011100101010011", 3872 => "1100111100111000", 3873 => "0010111011001000", 3874 => "1000010010101001", 3875 => "0000100001010100", 3876 => "1100111011110010", 3877 => "0111111101111101", 3878 => "1100111111111101", 3879 => "0010100110010000", 3880 => "0000001100101000", 3881 => "0001110111001000", 3882 => "0111000110010110", 3883 => "1111001011100110", 3884 => "1100100110010000", 3885 => "0101010100000010", 3886 => "0000000010010000", 3887 => "0100111001100110", 3888 => "0001101101100101", 3889 => "0011101110011000", 3890 => "0100101111110010", 3891 => "1100111001110011", 3892 => "0110001110110001", 3893 => "1000000001011111", 3894 => "1111111110100011", 3895 => "0001111011010011", 3896 => "0111110000111110", 3897 => "1100011011001001", 3898 => "0101001000110001", 3899 => "0001100100100110", 3900 => "1100011110100111", 3901 => "1101100010010001", 3902 => "1111100110011001", 3903 => "0111011100100101", 3904 => "0010110111110110", 3905 => "0111100111101000", 3906 => "0001001001101001", 3907 => "1101010010100001", 3908 => "0011001111010110", 3909 => "0001111111111010", 3910 => "1101000111010011", 3911 => "0110011011010000", 3912 => "1111000001100010", 3913 => "0101000100101111", 3914 => "0101101100101001", 3915 => "0010111100001100", 3916 => "1110010110100001", 3917 => "0100111010101100", 3918 => "0000110100110000", 3919 => "1111001111110101", 3920 => "0110100101001111", 3921 => "0111001010000010", 3922 => "0010000101110000", 3923 => "0111100101101010", 3924 => "1001000010100000", 3925 => "0010000100011010", 3926 => "0001001100110010", 3927 => "1111100000000110", 3928 => "0001111100001001", 3929 => "1010001011010000", 3930 => "1100001000010001", 3931 => "0100011000111101", 3932 => "0100000110100000", 3933 => "1100001100000110", 3934 => "1101110000000001", 3935 => "1100000011100101", 3936 => "0000011011011100", 3937 => "0010100100100011", 3938 => "0000011011000010", 3939 => "0001101111100000", 3940 => "1001111111010101", 3941 => "0011111100000010", 3942 => "0111010110010100", 3943 => "0101010111010000", 3944 => "1000010101110000", 3945 => "1010000010111111", 3946 => "1100001010010011", 3947 => "1001111010011111", 3948 => "0011100011101000", 3949 => "1000010000101000", 3950 => "1011010011001110", 3951 => "0010010111001001", 3952 => "0100110100011101", 3953 => "0101110011111011", 3954 => "1110001011101110", 3955 => "1001011001001000", 3956 => "0010000100001110", 3957 => "1100010110011110", 3958 => "1001101101000000", 3959 => "0010010000011011", 3960 => "0100001010001000", 3961 => "0100001111101000", 3962 => "1010011101100000", 3963 => "1011110110110000", 3964 => "0011101101110110", 3965 => "1001000000101101", 3966 => "1111110001000001", 3967 => "1010000000111101", 3968 => "1101110101110100", 3969 => "1001001000110001", 3970 => "0000101010110010", 3971 => "1010110011001001", 3972 => "0011101001001000", 3973 => "1110100011000110", 3974 => "1110000110100011", 3975 => "1100011110111111", 3976 => "1101000110101010", 3977 => "0100101001111101", 3978 => "0000011110110100", 3979 => "1001100110100011", 3980 => "1101000110110000", 3981 => "1110000100111110", 3982 => "1010010000000000", 3983 => "1111110000110110", 3984 => "0101010111010110", 3985 => "0011111011011000", 3986 => "0101011111110110", 3987 => "0000100001100001", 3988 => "0101001111000010", 3989 => "1100011111000001", 3990 => "1110001110101100", 3991 => "0010011000000110", 3992 => "0011000101111110", 3993 => "0010010101110010", 3994 => "1001111101110000", 3995 => "1111110101001101", 3996 => "0000010100001001", 3997 => "1101011110100101", 3998 => "0010110001010111", 3999 => "1001010110000000", 4000 => "1100110010110001", 4001 => "0011111111011001", 4002 => "1011000101110111", 4003 => "1010110010000101", 4004 => "1000110110110010", 4005 => "1001110010101101", 4006 => "0010000000011101", 4007 => "1011000000111011", 4008 => "1000010101011010", 4009 => "0010001000010100", 4010 => "1001011111110011", 4011 => "1001001011000010", 4012 => "1000111110011011", 4013 => "1011001110010000", 4014 => "0010000100010011", 4015 => "1111111110110101", 4016 => "0100111111110110", 4017 => "1001100010001111", 4018 => "1001010111110000", 4019 => "1011001000100001", 4020 => "1100000011001110", 4021 => "0010110001010100", 4022 => "0111101110111101", 4023 => "0110011110101100", 4024 => "0001001111011010", 4025 => "1110010011111001", 4026 => "1010000110111001", 4027 => "1101111110110101", 4028 => "1101110110110010", 4029 => "1011101011101010", 4030 => "1001111000100100", 4031 => "1001100110001100", 4032 => "1011001101111111", 4033 => "0000111001011101", 4034 => "1111111100011000", 4035 => "0111101110001100", 4036 => "1111001010001000", 4037 => "0110001111001001", 4038 => "1111010000110011", 4039 => "0101001111011001", 4040 => "1111100001001100", 4041 => "1011010000110000", 4042 => "0101001011000011", 4043 => "1110001001100110", 4044 => "0001001000100010", 4045 => "0010100000100110", 4046 => "1000011100001001", 4047 => "1010110111110011", 4048 => "1011010010111010", 4049 => "0011010000110000", 4050 => "0000111000111111", 4051 => "0111111001001000", 4052 => "1111100111000100", 4053 => "0110000011010100", 4054 => "0100011111101101", 4055 => "1110010010110010", 4056 => "1110110110010010", 4057 => "1011011100100111", 4058 => "1011011010101110", 4059 => "0100000001110111", 4060 => "1100111011101010", 4061 => "1010111111011110", 4062 => "0110010000000001", 4063 => "1110110000001101", 4064 => "0000001001101110", 4065 => "1001110000101110", 4066 => "1011010100011001", 4067 => "1110011011111010", 4068 => "0100110000110100", 4069 => "0101110001111100", 4070 => "0011110001010101", 4071 => "1101101001011001", 4072 => "0101110111111100", 4073 => "0010011011111000", 4074 => "1111100010000010", 4075 => "1111110011101011", 4076 => "1111111101110101", 4077 => "1001011100001010", 4078 => "1111110010110011", 4079 => "1011011001000100", 4080 => "0100010000010100", 4081 => "0100110110001101", 4082 => "0011110000101011", 4083 => "1101110001010011", 4084 => "0010110100110000", 4085 => "1100011110000001", 4086 => "0010101111110110", 4087 => "1000010011001000", 4088 => "1111111000011000", 4089 => "1010100101011000", 4090 => "0100101001011111", 4091 => "1101101110111111", 4092 => "1001111110001011", 4093 => "1100000011101001", 4094 => "0101010101110100", 4095 => "0110000010100010", 4096 => "0110011100011011", 4097 => "0010111101111100", 4098 => "1110000000001101", 4099 => "0010100101111110", 4100 => "1111000110110010", 4101 => "0100001001101100", 4102 => "1011001110101001", 4103 => "0101011011100100", 4104 => "0100101001010011", 4105 => "1011101011110111", 4106 => "0010100111010010", 4107 => "0011111101011011", 4108 => "0110001111011011", 4109 => "1110101001010101", 4110 => "1101111011100000", 4111 => "0100011011010111", 4112 => "1001110101011000", 4113 => "1000101110000001", 4114 => "0000110110100100", 4115 => "0111000100110011", 4116 => "1000011010111010", 4117 => "0100100110010000", 4118 => "0001001001111100", 4119 => "0100000011100111", 4120 => "1101001000001101", 4121 => "1011101111011010", 4122 => "0011000111111111", 4123 => "0111011100000000", 4124 => "1000011111001110", 4125 => "1000000001100101", 4126 => "0111100100010100", 4127 => "1101100000000010", 4128 => "1110111100100010", 4129 => "1000101100011110", 4130 => "0001001110100000", 4131 => "1001000101101100", 4132 => "1100011101100110", 4133 => "0100010110110110", 4134 => "0101010000000100", 4135 => "1000111101101001", 4136 => "1011000110011100", 4137 => "0000101011101110", 4138 => "1001100100101110", 4139 => "0000111101001000", 4140 => "1100101010111110", 4141 => "0111010111011100", 4142 => "1111011111111110", 4143 => "0010000111110000", 4144 => "0101111110110000", 4145 => "1111000011000100", 4146 => "1010111111000010", 4147 => "0100001101000101", 4148 => "1001010010100000", 4149 => "0110000010100110", 4150 => "0100110011011110", 4151 => "1101111000100011", 4152 => "1110100000100000", 4153 => "0011011011101101", 4154 => "1111011110101011", 4155 => "1001110001111100", 4156 => "1110010111100101", 4157 => "0101000111101000", 4158 => "1111010100001111", 4159 => "1000100100000101", 4160 => "1110000101010001", 4161 => "0111000010110001", 4162 => "1001111011110001", 4163 => "0000011010100000", 4164 => "1101110000101101", 4165 => "0010000011100010", 4166 => "1101110110001110", 4167 => "1001101101011000", 4168 => "1111000001010111", 4169 => "0010111001010001", 4170 => "1011110100010110", 4171 => "0001010111010110", 4172 => "0101000111110001", 4173 => "0010000110100000", 4174 => "0110111000001010", 4175 => "1110000110001100", 4176 => "1010101101011101", 4177 => "0101000011100010", 4178 => "0110010010111000", 4179 => "1101101110010111", 4180 => "0011000001011111", 4181 => "1111111110001111", 4182 => "0000000001100110", 4183 => "0111000110110011", 4184 => "0010110110010110", 4185 => "0010101000111110", 4186 => "1100110110100011", 4187 => "1001011001111101", 4188 => "1100111001011111", 4189 => "0110000010001001", 4190 => "0110110001110111", 4191 => "1001100001000011", 4192 => "1011100011010101", 4193 => "1000110110010011", 4194 => "1001110111101111", 4195 => "0010000100000011", 4196 => "0011101000111110", 4197 => "0100100100001110", 4198 => "0001011001001001", 4199 => "0011111111111111", 4200 => "0001111110000010", 4201 => "0000010110010101", 4202 => "0010111100100010", 4203 => "0111111100010001", 4204 => "0001110111100001", 4205 => "0011100000110110", 4206 => "0101100111110111", 4207 => "1010011110100010", 4208 => "1111111101100110", 4209 => "1010011111110001", 4210 => "1000011100110101", 4211 => "1100011001110101", 4212 => "1000101101001011", 4213 => "0101100000100010", 4214 => "0001110111100011", 4215 => "0100101100000100", 4216 => "0011001010000000", 4217 => "0111010111001100", 4218 => "0101000110100000", 4219 => "0011101100000111", 4220 => "0100101010000010", 4221 => "1101101001110110", 4222 => "0010111011011011", 4223 => "1110110111101101", 4224 => "1101011110111110", 4225 => "0111011010100010", 4226 => "0000011110101001", 4227 => "1101011010111100", 4228 => "0111011101001000", 4229 => "1000110111111000", 4230 => "0011101000010011", 4231 => "0111010001101111", 4232 => "0000001110110111", 4233 => "0000111110110001", 4234 => "1110000001100011", 4235 => "0110110111011101", 4236 => "0011111101001110", 4237 => "1100000010010000", 4238 => "0010110000110111", 4239 => "1111011000110111", 4240 => "0011110011110100", 4241 => "0001100111111001", 4242 => "1010001000010111", 4243 => "1000100111100011", 4244 => "0001100000001000", 4245 => "1011011011000101", 4246 => "1000001010111110", 4247 => "1010000011010000", 4248 => "1000100111000100", 4249 => "1101001101011101", 4250 => "1000111001001000", 4251 => "1101011011101111", 4252 => "0110100001100000", 4253 => "1010100111111011", 4254 => "0010100110100000", 4255 => "0101001001111011", 4256 => "1001000100111010", 4257 => "0111111011000111", 4258 => "0111110110101111", 4259 => "0101011101111011", 4260 => "1011101010110101", 4261 => "1001111111110010", 4262 => "1111111110110110", 4263 => "1100101000100000", 4264 => "1001011110000111", 4265 => "1101111111111110", 4266 => "0101101100100010", 4267 => "0010101110010010", 4268 => "1100100101001110", 4269 => "1100101111000010", 4270 => "1011101010110001", 4271 => "0010100010110001", 4272 => "0110101100110101", 4273 => "0110110110101111", 4274 => "1000000101001100", 4275 => "0000111100010000", 4276 => "0100101111100000", 4277 => "0001011110100100", 4278 => "0000101101111100", 4279 => "0010100100110101", 4280 => "1110001111111110", 4281 => "0100111001101010", 4282 => "1010010101011111", 4283 => "1001111111001011", 4284 => "1111001011000100", 4285 => "0110010011011100", 4286 => "0110011000111010", 4287 => "0111010101010110", 4288 => "1000101101101001", 4289 => "0100110100111100", 4290 => "0110110001010010", 4291 => "0100011010101000", 4292 => "0001100011001011", 4293 => "1000101101100100", 4294 => "1000010011111101", 4295 => "1010111110101100", 4296 => "0001100111101100", 4297 => "0010010001011011", 4298 => "1101110100011000", 4299 => "1111111110110111", 4300 => "0001000001100000", 4301 => "0001001110010111", 4302 => "0100001010011110", 4303 => "0111000010100001", 4304 => "0100101001100010", 4305 => "0111101001101101", 4306 => "0111001100100001", 4307 => "0001000010111101", 4308 => "1011011110110000", 4309 => "0011010100010111", 4310 => "0011011101011110", 4311 => "1011100001010100", 4312 => "0010110101100010", 4313 => "0111111110101100", 4314 => "1010100001110010", 4315 => "0001110110101010", 4316 => "0100110001101110", 4317 => "0110011101001000", 4318 => "1110101110011001", 4319 => "0101000110000110", 4320 => "0111001111001100", 4321 => "1101010101010011", 4322 => "1010000000000110", 4323 => "0001111010001101", 4324 => "1100001011100100", 4325 => "1100011100010100", 4326 => "0111100011101101", 4327 => "1110100110110100", 4328 => "1001111011011010", 4329 => "1001000001010011", 4330 => "1011011011101000", 4331 => "1011000101000100", 4332 => "1100111010110110", 4333 => "0011001000101111", 4334 => "1101111000110000", 4335 => "0011000111111110", 4336 => "0101011001101000", 4337 => "0001001000111101", 4338 => "1010010000010010", 4339 => "0001110111110100", 4340 => "1110100111101100", 4341 => "0111110100110110", 4342 => "1101110010111100", 4343 => "1101111011110010", 4344 => "0000101111001110", 4345 => "1011001001101101", 4346 => "0100110110011101", 4347 => "1111011100100110", 4348 => "0000000010000101", 4349 => "1100110101110100", 4350 => "0011110010001100", 4351 => "0111010101011101", 4352 => "0101100111000111", 4353 => "1101001100010110", 4354 => "1001101011001100", 4355 => "1000111000111110", 4356 => "1101000011111010", 4357 => "0110011110111101", 4358 => "0110011111011011", 4359 => "1000001001111101", 4360 => "1110001010100111", 4361 => "1011111101000101", 4362 => "1011000111111110", 4363 => "1111001111010001", 4364 => "1100000001010010", 4365 => "0101101010111001", 4366 => "0010110000110111", 4367 => "0100000010110001", 4368 => "1111000001100011", 4369 => "0001000000000011", 4370 => "1110000011010010", 4371 => "1110100000101010", 4372 => "1001011101100010", 4373 => "0010100011101100", 4374 => "0011001110100000", 4375 => "0010111000111010", 4376 => "1000111100001110", 4377 => "0100101101000011", 4378 => "0100101100100110", 4379 => "1100011000001111", 4380 => "0010011010101101", 4381 => "1100110111101111", 4382 => "0100000001111011", 4383 => "0101101001001011", 4384 => "0001010100110101", 4385 => "1011010011100010", 4386 => "1000100110010011", 4387 => "0111000110000011", 4388 => "1010001110000111", 4389 => "1111010110101100", 4390 => "1001001000110111", 4391 => "1010010000110101", 4392 => "1111011010100001", 4393 => "1100110111011000", 4394 => "0011011000000011", 4395 => "1111000101001011", 4396 => "0001000001100010", 4397 => "1010011010010100", 4398 => "1000001111110110", 4399 => "0110101101011000", 4400 => "1011110010011110", 4401 => "1000111001110010", 4402 => "1011010001101110", 4403 => "0011101101110110", 4404 => "0101010110110111", 4405 => "0111010101000100", 4406 => "1011100100000111", 4407 => "0111101000101011", 4408 => "0111010111010110", 4409 => "1000011101101100", 4410 => "0000010001011011", 4411 => "0011010101001000", 4412 => "0101110000101101", 4413 => "0000111001101011", 4414 => "0100010010111000", 4415 => "1100111110000010", 4416 => "0101001010001100", 4417 => "1110111111111111", 4418 => "1000000001011010", 4419 => "1101111110110111", 4420 => "0111000001100010", 4421 => "0101100100110110", 4422 => "0001101001110010", 4423 => "0000111110111010", 4424 => "1110110001001001", 4425 => "0001011100001101", 4426 => "1011111011110010", 4427 => "0001101110110100", 4428 => "1111000010101011", 4429 => "1000001000110110", 4430 => "1100000000011011", 4431 => "0111111001110111", 4432 => "1001011110011010", 4433 => "0111010001010010", 4434 => "0011000010111111", 4435 => "1101001111100000", 4436 => "1100100010001100", 4437 => "0001101110001100", 4438 => "1110011000100011", 4439 => "1011000110000111", 4440 => "0010101100000011", 4441 => "0000000010000101", 4442 => "1010100111001011", 4443 => "1011101101011110", 4444 => "0010110111111111", 4445 => "1000110101101001", 4446 => "0110100100100110", 4447 => "0111001111011000", 4448 => "1001010010001000", 4449 => "1100110111100101", 4450 => "0010010001000100", 4451 => "1100001011111000", 4452 => "1011001000110000", 4453 => "0011101001111010", 4454 => "1000110101101010", 4455 => "0011011111000010", 4456 => "0001010000000110", 4457 => "1010110011011010", 4458 => "1111000011110110", 4459 => "0110101101000110", 4460 => "1111111000100010", 4461 => "0010001011000001", 4462 => "1111111011010111", 4463 => "1010110011100111", 4464 => "1000001001011011", 4465 => "0001001101101100", 4466 => "0100111000100010", 4467 => "0100000110100001", 4468 => "0101000110000110", 4469 => "0001000100001001", 4470 => "0001100010001111", 4471 => "0111111000010000", 4472 => "1011000110010110", 4473 => "1110110110001011", 4474 => "0101110100000011", 4475 => "1100111101011110", 4476 => "1001001001010101", 4477 => "0111001110101110", 4478 => "0000111101001100", 4479 => "0010101000100000", 4480 => "1001110110101100", 4481 => "1011110111010101", 4482 => "1101010111001111", 4483 => "0001110011111011", 4484 => "0101011100011111", 4485 => "1101101001001100", 4486 => "0111111011001000", 4487 => "0111010001001110", 4488 => "1000000001100100", 4489 => "1111100100110101", 4490 => "0010011000000000", 4491 => "0100101110111010", 4492 => "1000001110100100", 4493 => "0011110001011001", 4494 => "0110011100100110", 4495 => "0111101011000111", 4496 => "1011111100110111", 4497 => "0001001110000110", 4498 => "0010001000100000", 4499 => "1010010011101110", 4500 => "1001001111001100", 4501 => "0110001011010111", 4502 => "0100100000001110", 4503 => "0000010010001011", 4504 => "0011000001010001", 4505 => "1111010000011101", 4506 => "0110110001000101", 4507 => "1000110000011111", 4508 => "0000100011110000", 4509 => "0000101000010001", 4510 => "1010010000011001", 4511 => "0001011011111101", 4512 => "0100110011110111", 4513 => "1011001001000110", 4514 => "0101110011010101", 4515 => "0010110001101011", 4516 => "1010001100100111", 4517 => "1101010011110001", 4518 => "0011100100100110", 4519 => "0110110110000001", 4520 => "1010110110001001", 4521 => "1100101100000001", 4522 => "1110101011001001", 4523 => "0110011000101101", 4524 => "0010010100110011", 4525 => "0100110000111111", 4526 => "1100101100111011", 4527 => "1001010101100100", 4528 => "0110010010110111", 4529 => "1101110110111110", 4530 => "1000101001111100", 4531 => "0101000000101010", 4532 => "1011101010011101", 4533 => "0011011011010010", 4534 => "1111101010111000", 4535 => "1011111100101101", 4536 => "0111010000100110", 4537 => "0010100011000011", 4538 => "1101111100010101", 4539 => "1110001000011000", 4540 => "1110101000001100", 4541 => "1000001001011000", 4542 => "1011000001110000", 4543 => "0100100001000010", 4544 => "1100101101100000", 4545 => "0000000001010000", 4546 => "1011011100111011", 4547 => "0011011010010011", 4548 => "0101100010011110", 4549 => "0110010011010001", 4550 => "0110101100000011", 4551 => "0101011001011101", 4552 => "1101101100101100", 4553 => "1001000111100011", 4554 => "0000110110010100", 4555 => "1100010101110010", 4556 => "0100101000100000", 4557 => "1100000100011010", 4558 => "0100100000110001", 4559 => "0001000101000100", 4560 => "1110100101100000", 4561 => "1110000100000110", 4562 => "0110010100011101", 4563 => "1100111010010110", 4564 => "1110111111101001", 4565 => "1011110001110000", 4566 => "1001101100100110", 4567 => "1110011010100010", 4568 => "0011011011001110", 4569 => "0110100010110111", 4570 => "1101011111001001", 4571 => "0100010000000111", 4572 => "1111011101000000", 4573 => "1101011001101011", 4574 => "0100000100110010", 4575 => "0011000110100110", 4576 => "0001001101101011", 4577 => "0011011011000100", 4578 => "0000110100001011", 4579 => "0000010011111110", 4580 => "1111111010101110", 4581 => "0110011010110101", 4582 => "0000100101110111", 4583 => "1010101001101010", 4584 => "0000111011011001", 4585 => "1010001111101110", 4586 => "0100110100010100", 4587 => "0101100110101110", 4588 => "0011000101100000", 4589 => "1111101100110011", 4590 => "1101110011011100", 4591 => "1101111110000111", 4592 => "1000011110010101", 4593 => "0111001101100101", 4594 => "1000001100111000", 4595 => "0000100100011111", 4596 => "0101001000101111", 4597 => "1110001010100100", 4598 => "1111101011010001", 4599 => "0110010000000011", 4600 => "0100101101011111", 4601 => "1101010111011101", 4602 => "1110011011101101", 4603 => "0001111101111001", 4604 => "0000100000100101", 4605 => "1100100111101011", 4606 => "0100001010110000", 4607 => "1100000001011110", 4608 => "0101000110010001", 4609 => "0001010010000000", 4610 => "0100110010000100", 4611 => "1110110001110111", 4612 => "0111000011001010", 4613 => "0000110111000011", 4614 => "1111010110001011", 4615 => "1111000011011101", 4616 => "0110000110101010", 4617 => "0000110001001000", 4618 => "1011111011001110", 4619 => "0110100011100010", 4620 => "1011100010001001", 4621 => "1110110011011100", 4622 => "0111100111101110", 4623 => "0001011011010001", 4624 => "0110000011110011", 4625 => "1010010110011111", 4626 => "1101010010000001", 4627 => "0000001101011100", 4628 => "0001111111001101", 4629 => "1110101011101000", 4630 => "1111101111101000", 4631 => "1101011100111110", 4632 => "1010010001100101", 4633 => "0011110011000001", 4634 => "1100001001010100", 4635 => "1000010100101101", 4636 => "0111001010100001", 4637 => "1100110010110110", 4638 => "0101110011100000", 4639 => "0001000001100101", 4640 => "0111111100011010", 4641 => "0011011110111101", 4642 => "0111110101110011", 4643 => "0011111011100001", 4644 => "0100000101110000", 4645 => "1100110101011010", 4646 => "1011001101010111", 4647 => "0011010100010011", 4648 => "1111000010000111", 4649 => "1010011110101101", 4650 => "1111010110011011", 4651 => "1111100001011001", 4652 => "0101001100100010", 4653 => "1101000100100101", 4654 => "0011100000000011", 4655 => "1001010001011011", 4656 => "1101000011000101", 4657 => "0011001110010001", 4658 => "1110101001100110", 4659 => "1101110001100110", 4660 => "1001000001101110", 4661 => "1111111011100100", 4662 => "0001110000011101", 4663 => "1111110000110100", 4664 => "0010011011111101", 4665 => "1011010011110111", 4666 => "0011001011111101", 4667 => "0010010110111111", 4668 => "0001100110110111", 4669 => "0010010011111000", 4670 => "1101010000110001", 4671 => "1011000110000100", 4672 => "1010111011101111", 4673 => "1101011110110011", 4674 => "0000111100110100", 4675 => "0110110101100110", 4676 => "0001001101010010", 4677 => "1011101100001110", 4678 => "0000101011010001", 4679 => "1111011101110011", 4680 => "0010111111001010", 4681 => "1010110010100100", 4682 => "0110000001111001", 4683 => "0000000000111001", 4684 => "1010010000000000", 4685 => "0100100100101100", 4686 => "1100000101010101", 4687 => "0101111101011010", 4688 => "1110110110101101", 4689 => "1101111000011001", 4690 => "1000010000101111", 4691 => "1010100001000010", 4692 => "0001001111101011", 4693 => "0001000111110101", 4694 => "1110000010010110", 4695 => "0011000100011101", 4696 => "0011111000100000", 4697 => "1110010110010010", 4698 => "1110101010001111", 4699 => "0111001110111001", 4700 => "1010110000010011", 4701 => "1011001010100000", 4702 => "0000001100111101", 4703 => "1000111000011011", 4704 => "0010000011101111", 4705 => "0100010001001010", 4706 => "0110010001001100", 4707 => "0101101011101011", 4708 => "1000011010011011", 4709 => "1110101000010101", 4710 => "1110000010111010", 4711 => "1000101110100010", 4712 => "0101000000100011", 4713 => "1101111001111111", 4714 => "0101010011001011", 4715 => "0111100110001110", 4716 => "0000000011011111", 4717 => "1011010000001001", 4718 => "1111111100011010", 4719 => "0100010100001101", 4720 => "1101101001100010", 4721 => "0111001001101011", 4722 => "0111100100101001", 4723 => "0110000110011111", 4724 => "0110011011001110", 4725 => "0000011011111110", 4726 => "1111111000011101", 4727 => "0011111000110000", 4728 => "1011100011100100", 4729 => "0010111111011110", 4730 => "0111101101110010", 4731 => "0110110001010000", 4732 => "1011101001111111", 4733 => "0100111011010011", 4734 => "0110110100000110", 4735 => "0001101011100011", 4736 => "0000010111111101", 4737 => "1000011111100001", 4738 => "0101011001001110", 4739 => "1111110101011000", 4740 => "0001001001011001", 4741 => "1100001001010010", 4742 => "0001100011000000", 4743 => "1101101110001110", 4744 => "1101100101011000", 4745 => "1101010110100110", 4746 => "0110100011110001", 4747 => "1001101010101010", 4748 => "1001100000100110", 4749 => "1000110010010100", 4750 => "0101110110000100", 4751 => "1101101011011111", 4752 => "0011100000100011", 4753 => "0101110100010101", 4754 => "0001101010101111", 4755 => "1110000011111010", 4756 => "0011111100001000", 4757 => "0000101010010011", 4758 => "0100111100001111", 4759 => "0011101001010101", 4760 => "0000010010001100", 4761 => "1110011101111100", 4762 => "1000011101111010", 4763 => "1110010110000011", 4764 => "0110010011110000", 4765 => "1110110000010111", 4766 => "1001110111100010", 4767 => "0100100011011000", 4768 => "1010111011010111", 4769 => "0000101111010101", 4770 => "0010101100010100", 4771 => "1111101101011100", 4772 => "0001000111011110", 4773 => "0101000111111111", 4774 => "1111100001011000", 4775 => "0110111101111010", 4776 => "1100111110000111", 4777 => "0110110101110011", 4778 => "0010011000100001", 4779 => "1110100011110100", 4780 => "0110111011011011", 4781 => "0100001011111000", 4782 => "0001000000110011", 4783 => "1101011011000011", 4784 => "1100000111011100", 4785 => "1011000010110001", 4786 => "1000110100001100", 4787 => "0001111100001100", 4788 => "1001000010001110", 4789 => "0101110010100101", 4790 => "0000000101111111", 4791 => "0011000001100000", 4792 => "1011001100100101", 4793 => "0100001010101001", 4794 => "1001000110000010", 4795 => "0011001101110000", 4796 => "0010000000000000", 4797 => "0101011100100100", 4798 => "0111010111000101", 4799 => "1100000010010011", 4800 => "1010101011010001", 4801 => "0111001000111011", 4802 => "1110101010110011", 4803 => "0001011011101110", 4804 => "1110011111100101", 4805 => "1000111010000000", 4806 => "0010001000111100", 4807 => "0000101100010110", 4808 => "0000001111100101", 4809 => "0111011010111001", 4810 => "1110100010110000", 4811 => "1111011000010100", 4812 => "0000101001001010", 4813 => "1101110011000100", 4814 => "0010001000100000", 4815 => "1100110001001100", 4816 => "1110101010011011", 4817 => "1001010010100010", 4818 => "0111101011010111", 4819 => "0110001110100001", 4820 => "1100011111011011", 4821 => "1110010001010111", 4822 => "1000111111111011", 4823 => "0000000100100101", 4824 => "0001111111011100", 4825 => "1010111011001100", 4826 => "1011111010100001", 4827 => "1011111100110111", 4828 => "1001000101011000", 4829 => "1010011101101101", 4830 => "1010000000110001", 4831 => "0110001011101011", 4832 => "1011111100110000", 4833 => "0100100001001101", 4834 => "0010000101011110", 4835 => "1011101111111010", 4836 => "0100000000110011", 4837 => "0001010000101111", 4838 => "1110101011000011", 4839 => "0101010010000010", 4840 => "0001010101101101", 4841 => "1100000010111011", 4842 => "1100000011100100", 4843 => "1000111011010001", 4844 => "1011000000101101", 4845 => "0001000110101101", 4846 => "1100000110100010", 4847 => "0001100101110110", 4848 => "1011010100000011", 4849 => "1111101110001100", 4850 => "1000001101100110", 4851 => "1111101011010000", 4852 => "1011010010011100", 4853 => "0101101000110110", 4854 => "1000101010100110", 4855 => "1011000001001110", 4856 => "1111000110010110", 4857 => "1001011110100000", 4858 => "1110110000111111", 4859 => "1010100000011100", 4860 => "0111101011101101", 4861 => "1111111011100010", 4862 => "1111110100111100", 4863 => "0010110100100001", 4864 => "1110000111010011", 4865 => "0011111111111111", 4866 => "0110010111100101", 4867 => "1010100110001011", 4868 => "1111011101110011", 4869 => "1110110001011110", 4870 => "1000101101011100", 4871 => "1100110000101010", 4872 => "0011001011101101", 4873 => "1111000011111010", 4874 => "1100101000111000", 4875 => "0100011101100111", 4876 => "0101010010101100", 4877 => "0010100000010110", 4878 => "0000001001001111", 4879 => "1001111101000110", 4880 => "0101000100000101", 4881 => "1110001000100111", 4882 => "1001110110001110", 4883 => "0000110001000010", 4884 => "0110101101011111", 4885 => "0110111011100010", 4886 => "1100110010110000", 4887 => "1011011111000110", 4888 => "0110101010101001", 4889 => "1001110000001011", 4890 => "1000010111000100", 4891 => "0001001110110010", 4892 => "1101000000111011", 4893 => "1110111010000100", 4894 => "1101101111110110", 4895 => "1100000001010101", 4896 => "1000000010100001", 4897 => "0010111001110011", 4898 => "1110100010101000", 4899 => "0010111100110001", 4900 => "0000001001001100", 4901 => "1001000011100010", 4902 => "1011000001100100", 4903 => "0111011011011101", 4904 => "0011011000101111", 4905 => "0100111110010100", 4906 => "0010100000010100", 4907 => "0101110111111100", 4908 => "1001110001111000", 4909 => "0010101001001111", 4910 => "0011010110101001", 4911 => "0010010101010000", 4912 => "0110000001111101", 4913 => "1011100000100101", 4914 => "0010111001000110", 4915 => "0000111110110000", 4916 => "1011111001011011", 4917 => "1101101011111011", 4918 => "1101000010111000", 4919 => "0110100001110001", 4920 => "1001010011100011", 4921 => "0111100110001010", 4922 => "0100001110001111", 4923 => "1110111000101100", 4924 => "0110100010010011", 4925 => "0101110100011011", 4926 => "1001110011111011", 4927 => "0001111101100100", 4928 => "0000110100011001", 4929 => "0111000001101001", 4930 => "1111100011000110", 4931 => "1010100000011111", 4932 => "0001100000111001", 4933 => "0101010110111100", 4934 => "1101111100000101", 4935 => "1011101111010111", 4936 => "1011101111110010", 4937 => "0001000010101010", 4938 => "0001101110101001", 4939 => "0011111010001011", 4940 => "0111111011100111", 4941 => "1000110100101111", 4942 => "0110110001010011", 4943 => "0001000001010000", 4944 => "0010100101100001", 4945 => "0100101110011011", 4946 => "0101110110101100", 4947 => "0001100000001110", 4948 => "0100010000111011", 4949 => "0110110010001001", 4950 => "0111001101101100", 4951 => "1011111101100001", 4952 => "1111010101011110", 4953 => "1011000110100000", 4954 => "1100101010100100", 4955 => "1001011111101000", 4956 => "0001110010000101", 4957 => "1000010001100101", 4958 => "0101011100111100", 4959 => "1111001111100011", 4960 => "0100100101011110", 4961 => "0011000010011101", 4962 => "0101100111001101", 4963 => "1000000001111101", 4964 => "0000010010011101", 4965 => "0111111100011000", 4966 => "1010001011000011", 4967 => "1001000101100010", 4968 => "1011010101111010", 4969 => "1101111100010001", 4970 => "1101110111000110", 4971 => "1111100110001011", 4972 => "1110010011010000", 4973 => "1011101000111011", 4974 => "1001101110100010", 4975 => "1111101011101100", 4976 => "0011111001100101", 4977 => "0000000101101001", 4978 => "0010011001000111", 4979 => "1000000101001010", 4980 => "0011110110001001", 4981 => "0100100010010001", 4982 => "0100010111101110", 4983 => "0010111101111101", 4984 => "0110010001011100", 4985 => "0101111000100101", 4986 => "1101010110100100", 4987 => "0101000001101110", 4988 => "1011010100100101", 4989 => "0100001011010110", 4990 => "1000111001001110", 4991 => "1011101111100110", 4992 => "0101000000001100", 4993 => "0011111000001010", 4994 => "1110100001011101", 4995 => "0100111110111110", 4996 => "1110011000100100", 4997 => "0111100111110101", 4998 => "0000111100111110", 4999 => "0010100010110010", 5000 => "1100100011111000", 5001 => "1110011000010011", 5002 => "1011010101110100", 5003 => "1101111001010001", 5004 => "1101110101101100", 5005 => "1001110111111100", 5006 => "1100001111000101", 5007 => "0111100111010010", 5008 => "1111010110100110", 5009 => "0001000010110100", 5010 => "1011111010001110", 5011 => "0011110011000111", 5012 => "1111000001011000", 5013 => "0011011001111000", 5014 => "1000000001010000", 5015 => "1000100111101101", 5016 => "1011101001110111", 5017 => "0110000001000111", 5018 => "0101001100000111", 5019 => "1110000100101011", 5020 => "0111001101010111", 5021 => "0100100101001011", 5022 => "0000110010100010", 5023 => "1110110011110111", 5024 => "1111100111001001", 5025 => "1110000100000111", 5026 => "0101010111001000", 5027 => "0010000001110000", 5028 => "1010001100011100", 5029 => "1010010110110010", 5030 => "1011000111001111", 5031 => "0011111000110101", 5032 => "0001001101100010", 5033 => "1001100011011011", 5034 => "1011110010101110", 5035 => "0000111111010001", 5036 => "0010111011111100", 5037 => "0110000111001100", 5038 => "1011010010010000", 5039 => "0100101101111000", 5040 => "1100011100010001", 5041 => "1100010111001110", 5042 => "0000111000001101", 5043 => "1110001100011000", 5044 => "1101001110101010", 5045 => "0110011001100111", 5046 => "0111001101011011", 5047 => "0001110110100011", 5048 => "0010010010000101", 5049 => "1111101110100001", 5050 => "1000101000011000", 5051 => "1110110001111001", 5052 => "0000101111010111", 5053 => "0001101011101011", 5054 => "0011010001011110", 5055 => "0101100000010110", 5056 => "0000011101100010", 5057 => "1011111101000000", 5058 => "1011010111011100", 5059 => "0101110110001011", 5060 => "0101110110011110", 5061 => "0110001011011110", 5062 => "0110000000111011", 5063 => "0010100110010001", 5064 => "1011110001001101", 5065 => "1011100000011101", 5066 => "1111001100101010", 5067 => "1101000011101000", 5068 => "0001100100001110", 5069 => "0101011101000100", 5070 => "1001100110100100", 5071 => "1010010100010011", 5072 => "1111010100111100", 5073 => "1001101000111111", 5074 => "1011100010110100", 5075 => "0101101000111010", 5076 => "0000011001101010", 5077 => "0101111010110000", 5078 => "0100111100110100", 5079 => "1110010011011111", 5080 => "1010100011011010", 5081 => "0101101001010001", 5082 => "1101110101110100", 5083 => "0001011101110111", 5084 => "1010110101101111", 5085 => "0001111000110110", 5086 => "0100101110010110", 5087 => "0111100110101000", 5088 => "0000001011110110", 5089 => "0001001010100010", 5090 => "0010010001010001", 5091 => "0000111101001110", 5092 => "0011110111111010", 5093 => "1011111001111010", 5094 => "0110010111001011", 5095 => "1001111010010111", 5096 => "0100010101111100", 5097 => "1001010111110100", 5098 => "1111101001011011", 5099 => "1111010101000101", 5100 => "1001011111101010", 5101 => "1111000000111111", 5102 => "1110110101000101", 5103 => "0010011000010111", 5104 => "1011101101000001", 5105 => "1000100100001100", 5106 => "1111010110001000", 5107 => "1000001110110111", 5108 => "1010100110011100", 5109 => "1000111101100110", 5110 => "0110111000000001", 5111 => "1100011101000100", 5112 => "1011000000100000", 5113 => "1000011010100101", 5114 => "0001011111000110", 5115 => "1010011111111000", 5116 => "0000111001000100", 5117 => "0011010100011010", 5118 => "0010001001011000", 5119 => "1111000110100000", 5120 => "1001000000000100", 5121 => "0110111101101000", 5122 => "0001011000110100", 5123 => "0110110100010010", 5124 => "0000000010011100", 5125 => "1011110101000110", 5126 => "1110000001010110", 5127 => "1001011111110000", 5128 => "1111011101111111", 5129 => "0000111011000101", 5130 => "1011111001011000", 5131 => "0011111000110001", 5132 => "0011010010011000", 5133 => "0110111100011100", 5134 => "1000101011111110", 5135 => "0000011111001100", 5136 => "1011011011110111", 5137 => "0001011011000110", 5138 => "0010101111101110", 5139 => "1110011110000011", 5140 => "0011110101001001", 5141 => "1001010100110110", 5142 => "0000000101100101", 5143 => "0000100101001110", 5144 => "1110010111111010", 5145 => "1011110001100001", 5146 => "0000001010111001", 5147 => "0101000000000110", 5148 => "1001111111001110", 5149 => "0010100111100110", 5150 => "1010101010110100", 5151 => "0100100111111100", 5152 => "0011100100011100", 5153 => "1010101011111001", 5154 => "0000000010110011", 5155 => "1011010000010001", 5156 => "1010011111000011", 5157 => "1101001101101111", 5158 => "0101011111000101", 5159 => "1011101111111000", 5160 => "1101100111000001", 5161 => "1011000111101001", 5162 => "0101110010010100", 5163 => "0010001010110000", 5164 => "1101101101011010", 5165 => "1001011111011001", 5166 => "0100010101010011", 5167 => "1000111010011101", 5168 => "0110110100001101", 5169 => "1110001111000011", 5170 => "1110110010101100", 5171 => "1110101101101100", 5172 => "0111000100101001", 5173 => "1001001100101101", 5174 => "1001111111010000", 5175 => "1110010110111110", 5176 => "1111000001110111", 5177 => "0001010100010010", 5178 => "1010110100100101", 5179 => "1101010100111100", 5180 => "1101000111000100", 5181 => "0010011110010010", 5182 => "0111111101111010", 5183 => "1100010010110010", 5184 => "0000001011101000", 5185 => "0100111000001010", 5186 => "1110001100100010", 5187 => "0111100101101100", 5188 => "0101011101011001", 5189 => "0101010011110001", 5190 => "0000110000101111", 5191 => "1110101110100100", 5192 => "1100110111011000", 5193 => "0001110110101001", 5194 => "0010010101111111", 5195 => "1110010011011101", 5196 => "0011010001010110", 5197 => "1110001100101101", 5198 => "0110110111111110", 5199 => "1001011000000000", 5200 => "0010101010010000", 5201 => "1110000101100101", 5202 => "0110010100101001", 5203 => "1010011111011101", 5204 => "0111000100000010", 5205 => "1010000100011100", 5206 => "0111010100100000", 5207 => "1010110011111111", 5208 => "0000000010110111", 5209 => "1100101001110111", 5210 => "1111010111011011", 5211 => "0101110000101010", 5212 => "1111110100000011", 5213 => "1010111110000011", 5214 => "0001110011001001", 5215 => "0010001000100101", 5216 => "1101100100100010", 5217 => "0111011000001001", 5218 => "0101011010110100", 5219 => "0011110101010001", 5220 => "0011111011101100", 5221 => "0111110101100001", 5222 => "1100001111100111", 5223 => "1100100001001001", 5224 => "0000011000000101", 5225 => "1110101001100110", 5226 => "1010110101101110", 5227 => "0010010000101101", 5228 => "0011010001101111", 5229 => "0000101101110100", 5230 => "0000101100110010", 5231 => "0110100110000101", 5232 => "1001001011110000", 5233 => "0000000000010110", 5234 => "1101111000010111", 5235 => "0111110111011101", 5236 => "1011100000110101", 5237 => "1000011100000110", 5238 => "1010110000010101", 5239 => "1110101100110011", 5240 => "0110011011010010", 5241 => "1011010100100000", 5242 => "0101100001111011", 5243 => "0110100011011101", 5244 => "0001000100111110", 5245 => "0011111010110101", 5246 => "0010001011101000", 5247 => "1101101001001000", 5248 => "0001110011101000", 5249 => "0100011000100001", 5250 => "0000111110001001", 5251 => "1011110101101010", 5252 => "1100111111011100", 5253 => "0010111011101010", 5254 => "0001001010111101", 5255 => "1111001010011011", 5256 => "1000110011011011", 5257 => "1101011111010010", 5258 => "0000001000000001", 5259 => "0101011100100100", 5260 => "1011111010000001", 5261 => "0111001001010010", 5262 => "0101110001010110", 5263 => "1001001010100000", 5264 => "1110010111110001", 5265 => "1111010111011011", 5266 => "1111001001110101", 5267 => "0001001110001100", 5268 => "1101111111011011", 5269 => "0000010101000100", 5270 => "0000110011101100", 5271 => "0010110001001110", 5272 => "0100101101010000", 5273 => "0111100010010101", 5274 => "1100111001001001", 5275 => "0100000011010010", 5276 => "0110001010101101", 5277 => "1000001011100010", 5278 => "1101000010011100", 5279 => "0000100111110111", 5280 => "0110010000010110", 5281 => "1010100001000101", 5282 => "0100001010001111", 5283 => "1010011011101010", 5284 => "1100000110001011", 5285 => "1000110000101101", 5286 => "1101001100000111", 5287 => "0101100101111100", 5288 => "1111011100011010", 5289 => "0011000100001001", 5290 => "1111011001010011", 5291 => "0010101010111111", 5292 => "0110101100110011", 5293 => "1111010101111000", 5294 => "1001001101000010", 5295 => "1001010111010001", 5296 => "1110100100000011", 5297 => "0011000101001001", 5298 => "1001010011110010", 5299 => "0011001100100111", 5300 => "1111101110010101", 5301 => "0011011011100010", 5302 => "1011001101100100", 5303 => "1011001111100100", 5304 => "0100110000001010", 5305 => "0010000000000000", 5306 => "0000111010110000", 5307 => "0101011111100100", 5308 => "0111101000000100", 5309 => "1100101001001101", 5310 => "0010110011110001", 5311 => "0100101011000110", 5312 => "0101101001110011", 5313 => "0101110110110001", 5314 => "0001011101111101", 5315 => "1010011110111101", 5316 => "0111001000010110", 5317 => "0001110110010011", 5318 => "1101101100110100", 5319 => "1111000110101010", 5320 => "1011110100011010", 5321 => "1100111000011110", 5322 => "0110111101000100", 5323 => "1010001101101000", 5324 => "1000101100100101", 5325 => "0011011100000101", 5326 => "0110111100101111", 5327 => "1100110101010011", 5328 => "0111111000101111", 5329 => "0110101000010001", 5330 => "0000111111010001", 5331 => "0101101010001101", 5332 => "1010110100010011", 5333 => "0100100101110000", 5334 => "0010000101101001", 5335 => "1110101100010010", 5336 => "0100100111000011", 5337 => "0001000011011000", 5338 => "0000110100111001", 5339 => "0001010010011101", 5340 => "1100101010101001", 5341 => "0110010101000101", 5342 => "0100110110110001", 5343 => "1101001101010011", 5344 => "0110001011010111", 5345 => "0010000111001010", 5346 => "1010111011001101", 5347 => "0111011010011111", 5348 => "1100011111011001", 5349 => "0111111010101110", 5350 => "1100101101111011", 5351 => "0111001110101010", 5352 => "1101010111000101", 5353 => "0100100000001110", 5354 => "1101100111101000", 5355 => "1001000010101100", 5356 => "1110000111101111", 5357 => "0100111010011110", 5358 => "1110110001101010", 5359 => "0001111100010000", 5360 => "1111101000100100", 5361 => "1101101110101010", 5362 => "0110010010100011", 5363 => "1110100000101001", 5364 => "1110110011101100", 5365 => "1101111000010100", 5366 => "1111110010000101", 5367 => "1011110001100000", 5368 => "1100101010001010", 5369 => "1110111011010101", 5370 => "0010000110000111", 5371 => "0010001000111111", 5372 => "0100110110101100", 5373 => "0100001010001111", 5374 => "1001101010100100", 5375 => "0010001111010010", 5376 => "0110110010100110", 5377 => "1011111000111110", 5378 => "1001101111111111", 5379 => "1111111011001101", 5380 => "0101100000100101", 5381 => "1000111011010011", 5382 => "0110011011100100", 5383 => "0110100011001101", 5384 => "1011101000000011", 5385 => "0000100101110110", 5386 => "1010001100000011", 5387 => "0111011001111100", 5388 => "1001010001001111", 5389 => "0110010001011100", 5390 => "0110110111001000", 5391 => "0011000101111010", 5392 => "1011010011011101", 5393 => "0111111101111010", 5394 => "1100111010100111", 5395 => "1110001110001011", 5396 => "1001001000000000", 5397 => "0101101111110100", 5398 => "1100100101011001", 5399 => "0101101101001101", 5400 => "0110111000011000", 5401 => "0100100111001111", 5402 => "1010010010101010", 5403 => "1000010100111011", 5404 => "1100100001001001", 5405 => "1111101100011111", 5406 => "1010010110111011", 5407 => "1100110010101010", 5408 => "1110100000101100", 5409 => "0110010110001011", 5410 => "1011101111100110", 5411 => "1010011100100101", 5412 => "1010110100011101", 5413 => "0000110111001111", 5414 => "0000101010011101", 5415 => "0101100110011101", 5416 => "0010101110000011", 5417 => "0110111110010100", 5418 => "0101010110011010", 5419 => "1111000101111011", 5420 => "1100010000110000", 5421 => "1101111101110000", 5422 => "0010111000110001", 5423 => "0001110011101001", 5424 => "0110110000011001", 5425 => "1010001001101110", 5426 => "1010101010010000", 5427 => "0011111110101100", 5428 => "0110001110100010", 5429 => "0010001010011011", 5430 => "0011110100111010", 5431 => "0101010010110100", 5432 => "0001110011001000", 5433 => "1001111011110101", 5434 => "0011111100001111", 5435 => "1001010011000101", 5436 => "1011000000100111", 5437 => "1010111011101010", 5438 => "1001111010011010", 5439 => "1000010011101111", 5440 => "0100100010111001", 5441 => "1100000011011000", 5442 => "0110110001111111", 5443 => "1010101111000101", 5444 => "0101110101000011", 5445 => "1011110100010010", 5446 => "0100011011000000", 5447 => "1100011000000010", 5448 => "0011000100011001", 5449 => "1100011101101000", 5450 => "0000011011010110", 5451 => "1101100110100111", 5452 => "0011000001110010", 5453 => "0101011101110101", 5454 => "1010110100001011", 5455 => "0010001110110011", 5456 => "0010011000100100", 5457 => "1010011100001101", 5458 => "1110011111111011", 5459 => "0011011110111100", 5460 => "1110110101100110", 5461 => "1010010001100001", 5462 => "0100111001110100", 5463 => "1100110011001001", 5464 => "0110110010100111", 5465 => "0111000001100001", 5466 => "1011011001000100", 5467 => "1111000111000011", 5468 => "1110110000000101", 5469 => "1010101011011100", 5470 => "1110001110011001", 5471 => "0110101011110000", 5472 => "1000101110011100", 5473 => "1110011110001001", 5474 => "0111011000110111", 5475 => "0001100000111011", 5476 => "0110001010010010", 5477 => "0110000001001100", 5478 => "1111111000011011", 5479 => "0001100000101101", 5480 => "1110011011101110", 5481 => "1110000100000111", 5482 => "0000111100011001", 5483 => "1101101100111110", 5484 => "1000110110001110", 5485 => "0100001001011010", 5486 => "1000011101111000", 5487 => "0000110011000101", 5488 => "0011110110001011", 5489 => "1111011110100000", 5490 => "0101000001111100", 5491 => "0000100110111111", 5492 => "1001101001001101", 5493 => "0010100001010101", 5494 => "0000110001111001", 5495 => "1101000110010111", 5496 => "0101011111111101", 5497 => "0010010110110101", 5498 => "1101010011010110", 5499 => "0111111010010001", 5500 => "1111111011000010", 5501 => "1101010000110011", 5502 => "1111110101110111", 5503 => "0010011101101011", 5504 => "1111110100110011", 5505 => "0111101111011000", 5506 => "0000011010110110", 5507 => "0101010111111110", 5508 => "1000110011001000", 5509 => "1101111111111001", 5510 => "1110111100011001", 5511 => "1001010000101010", 5512 => "0111001001101010", 5513 => "0000011111101100", 5514 => "1101010000101110", 5515 => "1111101101100111", 5516 => "0111001010001101", 5517 => "0000110110011010", 5518 => "1011101111110000", 5519 => "0101001001100001", 5520 => "1000110100101100", 5521 => "1100000010001000", 5522 => "0111101001011010", 5523 => "0000100011000101", 5524 => "1110101101100011", 5525 => "1001110110111000", 5526 => "0100000001101111", 5527 => "1001001111010110", 5528 => "0101100100111110", 5529 => "0000010001101111", 5530 => "0111011100110111", 5531 => "0100110111100100", 5532 => "0110101110010111", 5533 => "0010001101111111", 5534 => "0101110110100000", 5535 => "0001101000001111", 5536 => "0101011011111101", 5537 => "0110111001000001", 5538 => "0110101101000001", 5539 => "0001010010001111", 5540 => "1001011010110111", 5541 => "0110000111011111", 5542 => "0011111011110011", 5543 => "0100011111011101", 5544 => "0100110001001110", 5545 => "1010001110000010", 5546 => "0001101110111000", 5547 => "0001111111111000", 5548 => "0101111001010001", 5549 => "0011010010101111", 5550 => "1101010111010101", 5551 => "0101101000000011", 5552 => "1111011110010100", 5553 => "0010001001011011", 5554 => "1001001100001111", 5555 => "0110011111111100", 5556 => "0010001100101000", 5557 => "0101011011000111", 5558 => "1001011010100011", 5559 => "1100001001110001", 5560 => "0111001110011110", 5561 => "1011100100110000", 5562 => "1100001100101110", 5563 => "1100000110101010", 5564 => "1000000110111011", 5565 => "0110010101000110", 5566 => "0100000000010110", 5567 => "1001010011011111", 5568 => "0110111010110110", 5569 => "0011100001001101", 5570 => "0101010000011000", 5571 => "1011110110001011", 5572 => "0101011000001110", 5573 => "0001100000101001", 5574 => "0111011101000011", 5575 => "1101110101011011", 5576 => "1011110001111110", 5577 => "1100011111111011", 5578 => "0101110010101010", 5579 => "1111001001000101", 5580 => "1000001001000100", 5581 => "1001110110010001", 5582 => "0111000110001101", 5583 => "0111000000001101", 5584 => "1110011011101000", 5585 => "1001101001001100", 5586 => "1100010111101001", 5587 => "0010101001000010", 5588 => "0010110001011100", 5589 => "1110010111000101", 5590 => "1111011010011111", 5591 => "1101011110011101", 5592 => "1101000110101001", 5593 => "1110010010111001", 5594 => "1001100000101010", 5595 => "0101101110000110", 5596 => "1011001111110100", 5597 => "1010010101011011", 5598 => "0100001101100100", 5599 => "1111000100110111", 5600 => "1011100100111101", 5601 => "1000100010000100", 5602 => "1011110111010010", 5603 => "0000000000001110", 5604 => "0110010101000001", 5605 => "0010000111011011", 5606 => "0000001101001011", 5607 => "1001110000110110", 5608 => "0101001010110010", 5609 => "0000000001100001", 5610 => "1111010000110110", 5611 => "1010101111011000", 5612 => "0010111110101000", 5613 => "0101000011000111", 5614 => "0000001001011010", 5615 => "1011000001110010", 5616 => "0101101001101110", 5617 => "0000101011100100", 5618 => "1000101001010010", 5619 => "1010110100010001", 5620 => "0001110001011000", 5621 => "0111010000000100", 5622 => "1100101011000110", 5623 => "1111110000111110", 5624 => "0111001110010100", 5625 => "0011011000111110", 5626 => "1001011100001111", 5627 => "0000100111011001", 5628 => "1000111000011010", 5629 => "0001101000100111", 5630 => "0001111010010000", 5631 => "1111001010000111", 5632 => "0000111001110010", 5633 => "0101111100001000", 5634 => "0110101110101111", 5635 => "0111101101001101", 5636 => "0010001010000101", 5637 => "1101010001010100", 5638 => "0011100001111001", 5639 => "0101011111001110", 5640 => "1001110010010011", 5641 => "1101010110011110", 5642 => "1110101101011111", 5643 => "0110111110011100", 5644 => "1101001010000000", 5645 => "0100001100101110", 5646 => "1010000011000110", 5647 => "0100010010101110", 5648 => "1110000000100010", 5649 => "1101001000111010", 5650 => "0111110100111011", 5651 => "0000000010111011", 5652 => "0110111011001010", 5653 => "1010111000100110", 5654 => "0110100111110000", 5655 => "0110001111001101", 5656 => "1100000111011011", 5657 => "1011001101111010", 5658 => "0101011100001011", 5659 => "1111001011101010", 5660 => "1100011101010100", 5661 => "0011010011101100", 5662 => "1000011000010011", 5663 => "0111001010001010", 5664 => "0101010000000101", 5665 => "1100000010000001", 5666 => "1000010001100101", 5667 => "1000101000111100", 5668 => "1101010101101110", 5669 => "1011100011111110", 5670 => "0110010000011001", 5671 => "0000010000101011", 5672 => "0111011111111011", 5673 => "0111001010001001", 5674 => "1100111000011110", 5675 => "1001100001001001", 5676 => "0011110011100010", 5677 => "0010100010111010", 5678 => "0000100010111011", 5679 => "0101100110000110", 5680 => "0011111011001000", 5681 => "0110111000000101", 5682 => "1110011010011010", 5683 => "0101101100111011", 5684 => "1101100111101010", 5685 => "1101000000001100", 5686 => "1110011111010110", 5687 => "0001011001000010", 5688 => "0010011000101111", 5689 => "1101000111100010", 5690 => "0001110000110100", 5691 => "0010111010000110", 5692 => "1101111101100000", 5693 => "0010110111100010", 5694 => "1000001010010010", 5695 => "0111100000101011", 5696 => "0011111001010000", 5697 => "1010111111001110", 5698 => "1010000000011011", 5699 => "0000011101101110", 5700 => "0001000011101100", 5701 => "0110101111111011", 5702 => "1011111101110000", 5703 => "1111000111100011", 5704 => "1111010010111011", 5705 => "1100111010110101", 5706 => "0111111100001001", 5707 => "1111000011101001", 5708 => "0011100101100100", 5709 => "1110111101110000", 5710 => "1101010101011010", 5711 => "0111110000111010", 5712 => "1000100100101001", 5713 => "1000010000100110", 5714 => "1101101011010010", 5715 => "1101010110000110", 5716 => "1101011101011011", 5717 => "1011000011011000", 5718 => "0101101101000000", 5719 => "1111111101001001", 5720 => "0100001100111101", 5721 => "1001110010010001", 5722 => "0100011110010111", 5723 => "0110110101110000", 5724 => "1101011011100011", 5725 => "0100111011100000", 5726 => "0101111001110011", 5727 => "1001011000101010", 5728 => "1010000111010101", 5729 => "1000110001000111", 5730 => "1111001101011011", 5731 => "0110000101100001", 5732 => "0010100010011110", 5733 => "1101100110100110", 5734 => "0000001001100110", 5735 => "0110011010001001", 5736 => "0000100011001101", 5737 => "1101110101001011", 5738 => "0110111110000111", 5739 => "0100101001110111", 5740 => "0100110011001000", 5741 => "0100010000011011", 5742 => "0011101000111011", 5743 => "0010011001000100", 5744 => "0101000110001100", 5745 => "1110010010111011", 5746 => "0011110011010000", 5747 => "1010000100001010", 5748 => "1110100010011110", 5749 => "1011001010110100", 5750 => "0001001101001010", 5751 => "0001110101101011", 5752 => "0011101000110000", 5753 => "1000001101101011", 5754 => "1100101000011011", 5755 => "0010000001011010", 5756 => "1100010100000011", 5757 => "0100111110010011", 5758 => "1011010010001111", 5759 => "1011110111110100", 5760 => "0100000001110111", 5761 => "0000010101101010", 5762 => "0000011000110011", 5763 => "1010010001111000", 5764 => "0010100000000001", 5765 => "0100100101010111", 5766 => "1000011010001001", 5767 => "0100110011101000", 5768 => "0011111100100000", 5769 => "1011101101001111", 5770 => "1000110100110111", 5771 => "1111101000101000", 5772 => "0101111001001000", 5773 => "1111001100101101", 5774 => "1011011100110110", 5775 => "1011010110110100", 5776 => "0100010011101011", 5777 => "1000001111101000", 5778 => "1010010010101000", 5779 => "1001000000010111", 5780 => "1010100010001100", 5781 => "1001000110100100", 5782 => "0010100100000000", 5783 => "1111110111111011", 5784 => "1100000111011100", 5785 => "0100100000000001", 5786 => "0111110111011011", 5787 => "1001000101000001", 5788 => "0100110010000010", 5789 => "1011010100110110", 5790 => "0111010011101001", 5791 => "1110110001010001", 5792 => "0001100010001111", 5793 => "1000011110110111", 5794 => "0010011011100001", 5795 => "1011000101101001", 5796 => "0001010100001000", 5797 => "1000001100110011", 5798 => "1000100010110100", 5799 => "0001110101101001", 5800 => "1111000001000001", 5801 => "1111000111101010", 5802 => "1101000111110111", 5803 => "0110001011110111", 5804 => "0101100000110111", 5805 => "0101001001110011", 5806 => "0100001011011100", 5807 => "0001111010100010", 5808 => "0011011110000111", 5809 => "1001011001010001", 5810 => "0111110101100110", 5811 => "0101010001110111", 5812 => "1011011011010011", 5813 => "0010111000010010", 5814 => "0011010110011100", 5815 => "1110110010111000", 5816 => "0110110001101110", 5817 => "0110100011111001", 5818 => "0101111111000011", 5819 => "0100101010000011", 5820 => "1110011100110011", 5821 => "0000010001011100", 5822 => "1010110001100011", 5823 => "0111110001110000", 5824 => "1110011001010110", 5825 => "1001010000000110", 5826 => "0001001010010101", 5827 => "0111000101010110", 5828 => "1110101111111111", 5829 => "1101001010110000", 5830 => "0100100100000100", 5831 => "1010010001101001", 5832 => "1001111000101010", 5833 => "1010110010011010", 5834 => "1100011010110010", 5835 => "0111101110110011", 5836 => "0011110110100110", 5837 => "0001011111111011", 5838 => "0110011011010011", 5839 => "1110100001110000", 5840 => "0010111011101010", 5841 => "1100011010101111", 5842 => "0100000101111101", 5843 => "1100000001111001", 5844 => "1000000111110100", 5845 => "1101100101000000", 5846 => "0000111111001001", 5847 => "1101100000000000", 5848 => "1011001010110110", 5849 => "0100010011111010", 5850 => "1100010101000011", 5851 => "0111011111101000", 5852 => "0010100001111000", 5853 => "1001000001110111", 5854 => "0000100011001011", 5855 => "1001111011100110", 5856 => "0111110001111110", 5857 => "0111010101000000", 5858 => "1111011111101000", 5859 => "1011011000010100", 5860 => "0101011001001111", 5861 => "1111010101110000", 5862 => "0101011110101111", 5863 => "1111011010000001", 5864 => "0000110010100111", 5865 => "1000011001101100", 5866 => "1100001001110100", 5867 => "1010001101000000", 5868 => "1001010010011110", 5869 => "1100100000000100", 5870 => "0010100100101011", 5871 => "0100000100010001", 5872 => "1011010001011001", 5873 => "1110111000100001", 5874 => "0010101000011110", 5875 => "1010001101101100", 5876 => "1100110010011111", 5877 => "0101000010100100", 5878 => "0000010010001110", 5879 => "0001000110011010", 5880 => "0110011101101101", 5881 => "0001000100001110", 5882 => "0011101101011011", 5883 => "1001001011101000", 5884 => "0101111111111001", 5885 => "1001011001110110", 5886 => "0111001010011010", 5887 => "1100011000111010", 5888 => "1011111101101111", 5889 => "1011000110001101", 5890 => "1111011000110010", 5891 => "1010110101100100", 5892 => "1000111100001010", 5893 => "0010110110111000", 5894 => "1000011100110000", 5895 => "1000111111100011", 5896 => "0110000111100110", 5897 => "0001000011111000", 5898 => "1111010110010100", 5899 => "0110110000111001", 5900 => "0011011011011100", 5901 => "1010010001010001", 5902 => "0110100000001101", 5903 => "0101101001010010", 5904 => "1101111000100000", 5905 => "0110001101011011", 5906 => "1011011010111000", 5907 => "0110001110101111", 5908 => "0101110000100110", 5909 => "1110100111101000", 5910 => "1101011010101100", 5911 => "0011001010011000", 5912 => "0100001011100001", 5913 => "1100000000000111", 5914 => "0111010011011110", 5915 => "0001111001100011", 5916 => "0000000000010001", 5917 => "1111100100001010", 5918 => "1111110101100110", 5919 => "0110010011011100", 5920 => "1100100101010001", 5921 => "1110101010111011", 5922 => "1101001000011010", 5923 => "0100111100001000", 5924 => "0101111010010101", 5925 => "0100011100000101", 5926 => "0000111111110000", 5927 => "1100011010100010", 5928 => "1000101000011011", 5929 => "1011010010111101", 5930 => "0110101000101111", 5931 => "0100010001111010", 5932 => "0100101110110110", 5933 => "0011100010010011", 5934 => "0101000010111001", 5935 => "1010110101000100", 5936 => "1110100000101100", 5937 => "0000001000000101", 5938 => "0011110100111000", 5939 => "1001100101100001", 5940 => "1100001011010000", 5941 => "1110001111010110", 5942 => "0011100111000011", 5943 => "0110010101101001", 5944 => "1001101011000101", 5945 => "1101010011100111", 5946 => "0111101100001001", 5947 => "0001010000111001", 5948 => "1111111100101011", 5949 => "1110111110000001", 5950 => "0101101110011000", 5951 => "1001010111111100", 5952 => "1101110010100010", 5953 => "1111011100100010", 5954 => "1010010010100100", 5955 => "0101010000100101", 5956 => "0111011011001100", 5957 => "1100100000110001", 5958 => "1001000000110110", 5959 => "1000000101101001", 5960 => "0100110111000111", 5961 => "1100000010101100", 5962 => "1000110100010110", 5963 => "0011111010001001", 5964 => "1000010100100011", 5965 => "1111000101001101", 5966 => "1000101010111001", 5967 => "1101110000100001", 5968 => "0111100011010111", 5969 => "1101100101011010", 5970 => "0111010111101011", 5971 => "0111000111100001", 5972 => "1111010101010110", 5973 => "0011011101101011", 5974 => "1010111111001111", 5975 => "0000100010101010", 5976 => "1100111011100010", 5977 => "1110111110101010", 5978 => "1100111001000011", 5979 => "1001100101101000", 5980 => "0001001110111011", 5981 => "1010010010111010", 5982 => "0001000110010110", 5983 => "0111100011111111", 5984 => "0010100000000110", 5985 => "1010111001010110", 5986 => "1100101110011000", 5987 => "1111001011010000", 5988 => "0101100111101101", 5989 => "0000000100101110", 5990 => "1110000011001111", 5991 => "1100100001110101", 5992 => "0010111011111101", 5993 => "1111011001000111", 5994 => "1101001100110011", 5995 => "0011110111101111", 5996 => "1111100100110010", 5997 => "1111100010101011", 5998 => "0111100110010010", 5999 => "1010011001110001", 6000 => "1000110110010100", 6001 => "0011110111101011", 6002 => "1010001100110000", 6003 => "1110011000100011", 6004 => "1010111110110001", 6005 => "0011000100111110", 6006 => "0111011100110000", 6007 => "1101100101101100", 6008 => "0101011110101000", 6009 => "0101111010010110", 6010 => "0100110111000010", 6011 => "1111101100101110", 6012 => "1100011000011011", 6013 => "1100100110011111", 6014 => "0110111101010111", 6015 => "1000101010100010", 6016 => "1011010101111101", 6017 => "0010101011000101", 6018 => "1100000101111001", 6019 => "1110111010001110", 6020 => "0110011001111110", 6021 => "1011001000111010", 6022 => "0001010001000111", 6023 => "1100010100011001", 6024 => "1101010110101100", 6025 => "0100010111000100", 6026 => "0010111101010100", 6027 => "0111010010110111", 6028 => "1001111111011001", 6029 => "0110011000000011", 6030 => "1000110100001011", 6031 => "1001000001101001", 6032 => "0101011100001011", 6033 => "1101101010010101", 6034 => "0111000101101000", 6035 => "0011100100010010", 6036 => "0100000101100101", 6037 => "0101111000100010", 6038 => "0011011001111000", 6039 => "1010001011111100", 6040 => "1011100011001110", 6041 => "1011101010110011", 6042 => "1100001010100101", 6043 => "0110100010001101", 6044 => "1110011011001100", 6045 => "1011110111110100", 6046 => "1100000011001011", 6047 => "1110011111111100", 6048 => "1110001111110110", 6049 => "1101011110100000", 6050 => "0010010101110000", 6051 => "0100110011110010", 6052 => "0010011111010010", 6053 => "1001011110100011", 6054 => "0100001010111000", 6055 => "1110110101011000", 6056 => "1100011100011000", 6057 => "0110111010110111", 6058 => "1100000010011111", 6059 => "0100111100011101", 6060 => "1010011110111011", 6061 => "0000001101000110", 6062 => "0110011001101110", 6063 => "1011110001011001", 6064 => "0100000100011001", 6065 => "0000000001011100", 6066 => "1111010111111100", 6067 => "1011100101011100", 6068 => "0100001111001110", 6069 => "1101110100011011", 6070 => "0110001110001011", 6071 => "1100010110101101", 6072 => "1010111001010111", 6073 => "0011010111001000", 6074 => "0001111110010010", 6075 => "1011111001001111", 6076 => "0000011010110001", 6077 => "1100111010100011", 6078 => "0011010000111001", 6079 => "1010010101001000", 6080 => "1011111100101100", 6081 => "0110000011110101", 6082 => "1100100110111110", 6083 => "0100001100111011", 6084 => "0111101101111011", 6085 => "1010011100101010", 6086 => "0111010101010000", 6087 => "1011111000001101", 6088 => "1100011011110001", 6089 => "0110110001111001", 6090 => "0111111110000011", 6091 => "0100000001010001", 6092 => "1100010011100111", 6093 => "0100011010010111", 6094 => "1100111101100100", 6095 => "0111000101011101", 6096 => "1000111011010111", 6097 => "0001111101010110", 6098 => "1001011100110000", 6099 => "0010110000111100", 6100 => "1010010111111000", 6101 => "0111101101110010", 6102 => "1111110001011011", 6103 => "0101110011101011", 6104 => "1101110111001100", 6105 => "1000001100001100", 6106 => "0011011000000101", 6107 => "1111011000110001", 6108 => "1100011110010100", 6109 => "1001111001011110", 6110 => "0110010010111011", 6111 => "0110101010110111", 6112 => "1001111001101001", 6113 => "1000111000100001", 6114 => "1101101111110010", 6115 => "1001010010011100", 6116 => "0101010101111100", 6117 => "1101001110111101", 6118 => "1111111101100011", 6119 => "1011010111101001", 6120 => "0000100100101111", 6121 => "0001000011000100", 6122 => "0001110000001011", 6123 => "0000101001001001", 6124 => "1101101111101111", 6125 => "0100101000110000", 6126 => "1000001010011011", 6127 => "1011010110001011", 6128 => "0001001011010100", 6129 => "1010100011101010", 6130 => "0001011100111000", 6131 => "1101001011001100", 6132 => "1011101110111111", 6133 => "1011011101100000", 6134 => "1100001100101111", 6135 => "0101111110000011", 6136 => "0010110101111101", 6137 => "1100000011001001", 6138 => "1100110100011100", 6139 => "0110111011011000", 6140 => "1100011000011101", 6141 => "1011000110011101", 6142 => "0111000101000011", 6143 => "1011111000001011", 6144 => "1000100000110000", 6145 => "1010111101010111", 6146 => "0001010011010111", 6147 => "1011110101001111", 6148 => "1011011100000001", 6149 => "1010010011000101", 6150 => "0101111100100100", 6151 => "0011110001000100", 6152 => "0011101000111100", 6153 => "0101101111100001", 6154 => "0011101110100111", 6155 => "1111100111101010", 6156 => "0111000011011100", 6157 => "1000001001100000", 6158 => "1110110111000100", 6159 => "0000110110111000", 6160 => "0111111001100001", 6161 => "1000100011100011", 6162 => "1011110111001011", 6163 => "1011111001111101", 6164 => "1110011000111110", 6165 => "0100010011011111", 6166 => "1101101111001100", 6167 => "1010111011011001", 6168 => "0101111010110011", 6169 => "0011000010100100", 6170 => "1101010110001010", 6171 => "1111011001000110", 6172 => "1101001110010110", 6173 => "0000010010000110", 6174 => "0100101111001111", 6175 => "0101111001001100", 6176 => "1101000000111011", 6177 => "0111000010001111", 6178 => "1000010011110110", 6179 => "0111101010111110", 6180 => "0100110110001001", 6181 => "1011010111101010", 6182 => "0000011100100111", 6183 => "1110001011101101", 6184 => "1101110000011001", 6185 => "0101011111111100", 6186 => "0110000011000000", 6187 => "1111000001111010", 6188 => "1101000000100110", 6189 => "0111101101100100", 6190 => "1010111010010000", 6191 => "0011100000001000", 6192 => "1110100110111010", 6193 => "1010001110000110", 6194 => "1101110001101100", 6195 => "1011011011010001", 6196 => "1000001010100110", 6197 => "1110100100111010", 6198 => "0111011000000010", 6199 => "1011011101000110", 6200 => "1101110000101010", 6201 => "0100011111011011", 6202 => "1000101010101111", 6203 => "0111110100111001", 6204 => "0010000011100101", 6205 => "0010010011001101", 6206 => "0010111101100100", 6207 => "1101011011000011", 6208 => "0001011110011111", 6209 => "0000010010010011", 6210 => "1000111100000101", 6211 => "0111100010111000", 6212 => "1010110111011010", 6213 => "0010111000001001", 6214 => "1101111111100101", 6215 => "1111100111001101", 6216 => "0001110111011100", 6217 => "1001111111000001", 6218 => "0110001010001100", 6219 => "1101111011111011", 6220 => "1011101111110001", 6221 => "0000101111001111", 6222 => "0111011010011111", 6223 => "0011011000001000", 6224 => "0111100110011101", 6225 => "1010001011001101", 6226 => "1000101001110011", 6227 => "1110101000101010", 6228 => "0000010000111000", 6229 => "1010011000001011", 6230 => "1011000011100101", 6231 => "1110001110001111", 6232 => "1011111110011011", 6233 => "0001000111011110", 6234 => "0111111101010100", 6235 => "1101011100010101", 6236 => "0101100000000101", 6237 => "1110001010001111", 6238 => "1010011100000101", 6239 => "0000001100101101", 6240 => "1001111010010110", 6241 => "0101110101000111", 6242 => "1000110011010010", 6243 => "1101011111010100", 6244 => "0101101011101111", 6245 => "0111100001101010", 6246 => "1110001110000001", 6247 => "0000101000001001", 6248 => "1010110110100110", 6249 => "1111001000000001", 6250 => "1001011111000001", 6251 => "0011011100000111", 6252 => "0001111111001110", 6253 => "0101001110110011", 6254 => "1110110101011001", 6255 => "1010010000000000", 6256 => "1100101001110010", 6257 => "0101101010100001", 6258 => "1110111001011110", 6259 => "1011000100111001", 6260 => "1001111011010010", 6261 => "0010101100111101", 6262 => "0111111000000010", 6263 => "1101001111100111", 6264 => "1000010010000011", 6265 => "0110111000000101", 6266 => "1000111111010100", 6267 => "0100101001101110", 6268 => "1000011010101011", 6269 => "0111111110010110", 6270 => "0100111001100111", 6271 => "1111000101100011", 6272 => "0001011110110010", 6273 => "1110100011000001", 6274 => "1101101011101011", 6275 => "0010101111100001", 6276 => "0110110111111010", 6277 => "1010011011000011", 6278 => "1111000011001010", 6279 => "0000100101111010", 6280 => "1101101110111100", 6281 => "0101110110110101", 6282 => "1101100011100100", 6283 => "1101101000111011", 6284 => "0010101101100001", 6285 => "1110101111001110", 6286 => "1100111110111011", 6287 => "1101001111101110", 6288 => "0011001111000010", 6289 => "0011110111000001", 6290 => "1111010000101000", 6291 => "1001101000010101", 6292 => "1011110111011010", 6293 => "1011101000100011", 6294 => "1101110101000011", 6295 => "0100001110111100", 6296 => "0101001111011110", 6297 => "1001011110001111", 6298 => "0000101011100111", 6299 => "0011010101010100", 6300 => "0111111011010010", 6301 => "1111101010001011", 6302 => "0110100110110011", 6303 => "1001111110100011", 6304 => "0110000011010100", 6305 => "0001001111000101", 6306 => "1101110000011101", 6307 => "1000010010101111", 6308 => "0010111110101110", 6309 => "0010111111101110", 6310 => "0001010001011111", 6311 => "1010100010001111", 6312 => "1000010011001011", 6313 => "1101111101100010", 6314 => "1101111111100111", 6315 => "1011000100010011", 6316 => "1110000101010011", 6317 => "1101111001011001", 6318 => "1101101101110110", 6319 => "1100010010000110", 6320 => "1001010111110000", 6321 => "0101101111101100", 6322 => "0011001001110110", 6323 => "1000001100101000", 6324 => "0010111000000100", 6325 => "0100110000010111", 6326 => "1000110010111000", 6327 => "0001100011110100", 6328 => "0110011011000000", 6329 => "0001010000010001", 6330 => "0111100100101101", 6331 => "1000011011111111", 6332 => "1000000100001111", 6333 => "1110011000010111", 6334 => "1010100111111010", 6335 => "1100011000000101", 6336 => "1100011011000000", 6337 => "1111110001100011", 6338 => "1000000010100000", 6339 => "1001110100011111", 6340 => "1001101110001110", 6341 => "1100001110000111", 6342 => "0101000110111100", 6343 => "1000011011010101", 6344 => "0101101000100011", 6345 => "0111101011011010", 6346 => "0101010110110100", 6347 => "0100110011101010", 6348 => "1001111011111100", 6349 => "1101000100011110", 6350 => "1000100101110111", 6351 => "1010101110000101", 6352 => "1011001011000010", 6353 => "0000011001111110", 6354 => "1000101100001110", 6355 => "1010100111111110", 6356 => "0111110001011101", 6357 => "1011000011010001", 6358 => "0110110101100101", 6359 => "0110001000000110", 6360 => "1010000010101000", 6361 => "0111100101110001", 6362 => "1100100100001111", 6363 => "1000010111100111", 6364 => "0111100100111111", 6365 => "1101010100011000", 6366 => "0000111110001110", 6367 => "0010000101101001", 6368 => "0000010000110101", 6369 => "1011110010111010", 6370 => "0101011000111010", 6371 => "0111001000001110", 6372 => "0111010001010111", 6373 => "1110110110010011", 6374 => "0001100010010001", 6375 => "0011101100000000", 6376 => "1100000000101110", 6377 => "1010111000110100", 6378 => "1001010010111111", 6379 => "1110001101010110", 6380 => "1000100100100000", 6381 => "1111010000100011", 6382 => "0010100010101110", 6383 => "1010101010111101", 6384 => "1101100101001100", 6385 => "0110100000011010", 6386 => "1001001111010000", 6387 => "0111000000101001", 6388 => "0111111001101100", 6389 => "0100100010001000", 6390 => "1110001001111001", 6391 => "1001100011111110", 6392 => "1001001001001000", 6393 => "1010110101100001", 6394 => "1100110001111111", 6395 => "1010011010100111", 6396 => "0000010101011000", 6397 => "0110110100000101", 6398 => "1011011000001100", 6399 => "1011111000001101", 6400 => "0111101011100111", 6401 => "0111100100010100", 6402 => "1011000010111010", 6403 => "0011010100111110", 6404 => "0111000010111010", 6405 => "0010001110111111", 6406 => "0111101000001110", 6407 => "1110011001101001", 6408 => "1101101000111111", 6409 => "1000100011110011", 6410 => "1101000100010111", 6411 => "1110000011001100", 6412 => "0010011001100000", 6413 => "0100100101110111", 6414 => "1111011001011100", 6415 => "1101011101000100", 6416 => "1110111001101100", 6417 => "0011101111000110", 6418 => "1100111110001001", 6419 => "0100000100110100", 6420 => "1001101001110011", 6421 => "0010001001000110", 6422 => "0111001000100011", 6423 => "0011101111111101", 6424 => "1010011000000100", 6425 => "1010101001001011", 6426 => "0001111001100101", 6427 => "0100001110110110", 6428 => "0011001100011000", 6429 => "1110110100001100", 6430 => "0100100101011010", 6431 => "1100011001000111", 6432 => "1110110101001100", 6433 => "0111100111010111", 6434 => "0000010110110101", 6435 => "0011111010111001", 6436 => "0010011000111110", 6437 => "1101000011011101", 6438 => "0111101100001101", 6439 => "1101001100000111", 6440 => "0101100000100001", 6441 => "1110010101011001", 6442 => "1011101100010010", 6443 => "1110111000111101", 6444 => "1000100101100101", 6445 => "0011001111001011", 6446 => "0111001001001001", 6447 => "0011100000100010", 6448 => "1010011010000100", 6449 => "0011100001010101", 6450 => "1111010111100010", 6451 => "1110000001011011", 6452 => "0001011100011101", 6453 => "0110101110001111", 6454 => "0100011010100000", 6455 => "0110011000110000", 6456 => "0110000011100110", 6457 => "0010110000111111", 6458 => "0010110001011100", 6459 => "1010110110111001", 6460 => "0111111100110010", 6461 => "0100100010010101", 6462 => "0011111101001010", 6463 => "0110111101100100", 6464 => "1011011110100000", 6465 => "0011000000000010", 6466 => "1000111101110111", 6467 => "1011100010010111", 6468 => "0101111111111011", 6469 => "1111001000010000", 6470 => "0001100110010000", 6471 => "0011000101101000", 6472 => "0011010001000010", 6473 => "0101011111101011", 6474 => "0111101101100011", 6475 => "1001101010001101", 6476 => "1011001110001110", 6477 => "1001011010111001", 6478 => "1011000110111110", 6479 => "1001001100011111", 6480 => "1001000110011001", 6481 => "1100100100100111", 6482 => "0010010011111011", 6483 => "0010011000001111", 6484 => "1001001001010001", 6485 => "0010001100110101", 6486 => "0011101100111111", 6487 => "1000101101101010", 6488 => "1100010001010110", 6489 => "1101110101101011", 6490 => "1010100010111100", 6491 => "0111011000111111", 6492 => "1100010011100101", 6493 => "0101001000101000", 6494 => "0100001001011101", 6495 => "1100001101111000", 6496 => "1110100010110111", 6497 => "0110110011010100", 6498 => "1110101111010110", 6499 => "1110110001001011", 6500 => "0000100110100011", 6501 => "0101010001001101", 6502 => "1110110111111101", 6503 => "1010011001001111", 6504 => "0111101110111110", 6505 => "0000100111101001", 6506 => "0011110010111001", 6507 => "1100010100111111", 6508 => "1111111101011011", 6509 => "1101001010001110", 6510 => "1011100110000101", 6511 => "0000011101000101", 6512 => "1100010101001110", 6513 => "0000011010110010", 6514 => "0100010111100010", 6515 => "1000010101111100", 6516 => "1111111111101001", 6517 => "1100101101101100", 6518 => "1000001101110001", 6519 => "0010101000000000", 6520 => "0000010110000101", 6521 => "0001011111010000", 6522 => "1010001101101001", 6523 => "0100110011001010", 6524 => "1111001010000010", 6525 => "1110100101111111", 6526 => "0111111010010100", 6527 => "0111111100100101", 6528 => "1110011111111101", 6529 => "0000101111110000", 6530 => "1001111110001110", 6531 => "1011011011010101", 6532 => "1010011011100010", 6533 => "1101111100000010", 6534 => "1010111001110110", 6535 => "0100001001000010", 6536 => "0110111100110011", 6537 => "0111001011110001", 6538 => "0001010100010100", 6539 => "0000111000111100", 6540 => "1110101010110011", 6541 => "0010110101010110", 6542 => "0010100010100110", 6543 => "0110110011110111", 6544 => "1010111110111101", 6545 => "0100110100010111", 6546 => "0001011101001110", 6547 => "1101110110010010", 6548 => "0100110000110001", 6549 => "0101101011001111", 6550 => "1100100111100111", 6551 => "0101000110100110", 6552 => "1111110000010110", 6553 => "0001100001000110", 6554 => "0110011010010000", 6555 => "1111000011100100", 6556 => "0000100111001000", 6557 => "0111101110100000", 6558 => "0101100101101101", 6559 => "1010010000011010", 6560 => "1110000111001101", 6561 => "1001101111001001", 6562 => "0101101101101100", 6563 => "0111000001110000", 6564 => "1100010000011110", 6565 => "0111000000110000", 6566 => "0011000101101100", 6567 => "0101010100011001", 6568 => "1110100110000001", 6569 => "1011110111010000", 6570 => "1101101011011011", 6571 => "1010010110101111", 6572 => "0111010100111001", 6573 => "1101000110111000", 6574 => "0101110110111001", 6575 => "0111011010000000", 6576 => "1110101110100100", 6577 => "0000000000010000", 6578 => "0101011001101100", 6579 => "1101011010000001", 6580 => "0000001110011011", 6581 => "0010011111010111", 6582 => "1011010011011010", 6583 => "0110011001001110", 6584 => "1011100100101011", 6585 => "1001011000111010", 6586 => "1101100000111100", 6587 => "1100101000100010", 6588 => "1110101110000100", 6589 => "0011001011100001", 6590 => "0111101110100110", 6591 => "0111001011101101", 6592 => "1001001011000010", 6593 => "1101111000101011", 6594 => "0100101100101010", 6595 => "0000111110111110", 6596 => "1001111010000000", 6597 => "0101110000110000", 6598 => "0011011110100000", 6599 => "1000100001010001", 6600 => "0001011001001000", 6601 => "1010100001110011", 6602 => "0110111100101100", 6603 => "0101011111111000", 6604 => "1100100010001101", 6605 => "0001101010111110", 6606 => "1001111100010100", 6607 => "1100001000111111", 6608 => "1010111011010100", 6609 => "0001100110010001", 6610 => "0000110011011000", 6611 => "1110110111101100", 6612 => "1011011000010111", 6613 => "0000111100010110", 6614 => "0100100110011011", 6615 => "1000011010010001", 6616 => "0001110100111010", 6617 => "0011110001010001", 6618 => "1111010010001001", 6619 => "0001010110110010", 6620 => "0111001001110100", 6621 => "1000101011000011", 6622 => "0111101100000011", 6623 => "1000011010001101", 6624 => "0000100011000000", 6625 => "1010111001011111", 6626 => "1101100001111010", 6627 => "0100001001111001", 6628 => "1010100101000001", 6629 => "0100011111001010", 6630 => "0011001100000100", 6631 => "1011011111000001", 6632 => "0010100111010010", 6633 => "1110010001101011", 6634 => "0101111111000111", 6635 => "0111101000111001", 6636 => "1001011111110110", 6637 => "1001000001100100", 6638 => "0000000110010000", 6639 => "0011100001010001", 6640 => "0000110010001011", 6641 => "1000001000010101", 6642 => "1110010100010100", 6643 => "1111010100110100", 6644 => "0011101101111111", 6645 => "1011111000101011", 6646 => "1100011000011011", 6647 => "0101111010001011", 6648 => "1111010100111010", 6649 => "0111000110011010", 6650 => "0100110111001001", 6651 => "0100110100111100", 6652 => "1101100110110000", 6653 => "0001101010101110", 6654 => "1001010000111111", 6655 => "0111010100111100", 6656 => "1011100111000111", 6657 => "1001100101100110", 6658 => "0010110011100011", 6659 => "1011100001010111", 6660 => "1100001110000011", 6661 => "0010000111010100", 6662 => "0011000100010011", 6663 => "1000100010001011", 6664 => "0001011010011001", 6665 => "0001111111010101", 6666 => "1111100100101010", 6667 => "1110011000010000", 6668 => "1000110000111100", 6669 => "0110110000011110", 6670 => "1110011101110111", 6671 => "1111000010011100", 6672 => "0111101111100000", 6673 => "1001110010000011", 6674 => "1111110110111100", 6675 => "1010110101001111", 6676 => "0100001110001101", 6677 => "1100100110110000", 6678 => "1100011011100101", 6679 => "1001110101000010", 6680 => "0001001111000111", 6681 => "0000011000001001", 6682 => "1110001101111000", 6683 => "0101010000100110", 6684 => "0100101110001101", 6685 => "0100101100010100", 6686 => "1011010010111100", 6687 => "0010101110001001", 6688 => "0101011110010111", 6689 => "0010011011100110", 6690 => "1110100110100100", 6691 => "0111000111011100", 6692 => "0111110111111001", 6693 => "0111000011110001", 6694 => "1001001000010011", 6695 => "0010111101101110", 6696 => "1010010000101010", 6697 => "1000001111001000", 6698 => "0111010000110011", 6699 => "0000110100011101", 6700 => "1101100111010010", 6701 => "0001111110011111", 6702 => "1001000111110010", 6703 => "1000001000100100", 6704 => "1011100101010001", 6705 => "0111100101000101", 6706 => "1010011101011001", 6707 => "1100101001110010", 6708 => "0010000001000101", 6709 => "1100101101011001", 6710 => "1010011000000101", 6711 => "0010011000110000", 6712 => "0110110101000011", 6713 => "1101111101111010", 6714 => "0010111000011101", 6715 => "0101111001010111", 6716 => "0111000000001110", 6717 => "1000110101110001", 6718 => "0111000110001111", 6719 => "1110000010001100", 6720 => "0100110001111001", 6721 => "1010110101110101", 6722 => "0100101011001010", 6723 => "1111010001011111", 6724 => "0011100010110000", 6725 => "0011101000011011", 6726 => "1011011110101000", 6727 => "1101100001101010", 6728 => "0001100010010001", 6729 => "0001000110010111", 6730 => "1000011110000111", 6731 => "1011100001001100", 6732 => "1111111010001101", 6733 => "0110101111111100", 6734 => "0110001110001001", 6735 => "1101101001101101", 6736 => "0101011101111000", 6737 => "0000110101110101", 6738 => "1110111110111000", 6739 => "0001001010111010", 6740 => "0010011101100110", 6741 => "0110100011011111", 6742 => "0111010110110110", 6743 => "1000100110101010", 6744 => "0001111000111011", 6745 => "1101111000000010", 6746 => "1100000001010110", 6747 => "0001010101011111", 6748 => "1111011111110000", 6749 => "0010011000100101", 6750 => "0101110000010111", 6751 => "0111110111010101", 6752 => "1010101101110100", 6753 => "0110010011001100", 6754 => "1100100000000001", 6755 => "0100101010111110", 6756 => "0110011110111010", 6757 => "1000010010010110", 6758 => "1111000001101000", 6759 => "0011011100110011", 6760 => "1101110100001010", 6761 => "1100100110101011", 6762 => "0100111000110011", 6763 => "1010010100001111", 6764 => "0111000011010000", 6765 => "1101011010101000", 6766 => "1011110100101110", 6767 => "1111110010011010", 6768 => "0000001110111110", 6769 => "1001000111011011", 6770 => "1001100100110001", 6771 => "0000010110011001", 6772 => "1001110000001001", 6773 => "1101111110101011", 6774 => "0110101101010001", 6775 => "0100001101011000", 6776 => "0100001111101100", 6777 => "0101101110000100", 6778 => "1100000101010000", 6779 => "0101001001101001", 6780 => "1010000111111001", 6781 => "0100101010110100", 6782 => "0011110110010001", 6783 => "1000100100101010", 6784 => "1111101101110000", 6785 => "0100111001110101", 6786 => "0000110001000100", 6787 => "0101101100100110", 6788 => "0000001001100110", 6789 => "1101010010110111", 6790 => "0001011000101000", 6791 => "1111010111010001", 6792 => "1000001010101011", 6793 => "0100001010010010", 6794 => "1101010000011101", 6795 => "0111001000110101", 6796 => "0001000111000000", 6797 => "0001110100100101", 6798 => "1000000001001010", 6799 => "0011100110111001", 6800 => "1001000011101100", 6801 => "1010000010100000", 6802 => "0011001101100001", 6803 => "0101011100000100", 6804 => "1101101011111110", 6805 => "1000001010101110", 6806 => "0000010101111100", 6807 => "0101111010100110", 6808 => "0101100110001111", 6809 => "1110100000000001", 6810 => "0111000010100111", 6811 => "0110000011100111", 6812 => "0001101101111011", 6813 => "1110100110011010", 6814 => "0000010100111101", 6815 => "0110000010000000", 6816 => "0101010110100010", 6817 => "0110101000010001", 6818 => "1001101000101000", 6819 => "0101110110011110", 6820 => "1001100001011011", 6821 => "1000011011100101", 6822 => "1001011011101000", 6823 => "0011110000110111", 6824 => "0010000100110000", 6825 => "0100100101010101", 6826 => "1111001011000011", 6827 => "1010010111011110", 6828 => "0101110101011000", 6829 => "1010001101000110", 6830 => "0111001011001110", 6831 => "1000010000001010", 6832 => "1001101100100111", 6833 => "0100010111110111", 6834 => "0010011110001101", 6835 => "0111001010001101", 6836 => "0001011001010001", 6837 => "1101101000000011", 6838 => "0010100011010110", 6839 => "0101011000111101", 6840 => "0101000110001111", 6841 => "1011011110001100", 6842 => "1111001001010111", 6843 => "1110011100101100", 6844 => "0010101110011000", 6845 => "1101100110111100", 6846 => "0010000110101011", 6847 => "1001010000110110", 6848 => "1001011010001110", 6849 => "1011100000010110", 6850 => "0001010011010011", 6851 => "1011111110001111", 6852 => "0010001110100100", 6853 => "1000110010011001", 6854 => "0000111101111111", 6855 => "0101101010000011", 6856 => "1111100100000111", 6857 => "0011011110010011", 6858 => "0111100100101000", 6859 => "0011101001001110", 6860 => "0101110010000110", 6861 => "0001000110010101", 6862 => "0111101010000011", 6863 => "0000100011001100", 6864 => "1010110101111000", 6865 => "0110100010001011", 6866 => "1110010111111110", 6867 => "0011111101110011", 6868 => "0011111100100111", 6869 => "1001111011001110", 6870 => "1000000000101101", 6871 => "1111101001000000", 6872 => "0000111000110100", 6873 => "0111011101111010", 6874 => "0000010011110000", 6875 => "0000011100001011", 6876 => "1111110101001110", 6877 => "1010000001010101", 6878 => "1111100000000111", 6879 => "0101101101100010", 6880 => "1001100011000111", 6881 => "1101001011010100", 6882 => "0011100111000101", 6883 => "0101001101111011", 6884 => "1110001010111100", 6885 => "1010000010111100", 6886 => "1000110100101010", 6887 => "1010010111101101", 6888 => "0100000010011000", 6889 => "1000101110101111", 6890 => "0010010010100100", 6891 => "0111010001000100", 6892 => "1111010000010110", 6893 => "0000010011001111", 6894 => "1110101100110110", 6895 => "1001010000010010", 6896 => "1001110011001110", 6897 => "0011111100001011", 6898 => "0111011100000010", 6899 => "1100001011101101", 6900 => "0011001000001000", 6901 => "0010000101011100", 6902 => "0110101000011111", 6903 => "0000011101011011", 6904 => "1001001000101110", 6905 => "1100110000011111", 6906 => "1100011111010101", 6907 => "1000011010011110", 6908 => "1000011111011111", 6909 => "1000000010111111", 6910 => "0001110101111101", 6911 => "0111000111100111", 6912 => "1110110010000100", 6913 => "1011011100000110", 6914 => "1101010001010100", 6915 => "1101010110101010", 6916 => "0111001010111010", 6917 => "0010001000001000", 6918 => "1111000100111001", 6919 => "1101011011010010", 6920 => "0001001000111111", 6921 => "0111101000001100", 6922 => "0111100111000000", 6923 => "0001110100111101", 6924 => "0011111011110100", 6925 => "0000111110100101", 6926 => "1111111011001111", 6927 => "0110111011111011", 6928 => "0101000011100010", 6929 => "0110001100001110", 6930 => "1100111001011010", 6931 => "1001111001011011", 6932 => "0000001111111100", 6933 => "0101011010010000", 6934 => "0011100001100011", 6935 => "1010110111000101", 6936 => "1100100111011101", 6937 => "0000100110111010", 6938 => "0000001111001101", 6939 => "1101000111010011", 6940 => "1011011010110001", 6941 => "1110010101000111", 6942 => "1010101000111111", 6943 => "0010011111100001", 6944 => "0011110110111100", 6945 => "0111100100100010", 6946 => "1011100100110111", 6947 => "0111101110111010", 6948 => "1101001000100001", 6949 => "0101001001001001", 6950 => "1111111010111111", 6951 => "1010101001110001", 6952 => "1000001111011110", 6953 => "0000110101100101", 6954 => "1010110110011001", 6955 => "1100100100101011", 6956 => "1110111001011011", 6957 => "1011011001100111", 6958 => "1100010110011101", 6959 => "0110011001010100", 6960 => "0101001000111000", 6961 => "0001000011101111", 6962 => "1100110001100100", 6963 => "0100000101111010", 6964 => "1010001010101000", 6965 => "1001011100011000", 6966 => "0011111011001110", 6967 => "0101110101100011", 6968 => "1001110001000001", 6969 => "0010011111101110", 6970 => "0110111101101110", 6971 => "1101000101100111", 6972 => "1001101010010111", 6973 => "1100111000001011", 6974 => "0011100000110010", 6975 => "1011110100110111", 6976 => "0111110001101111", 6977 => "1000001001111000", 6978 => "1101111111010000", 6979 => "1100110001100000", 6980 => "1000010001111110", 6981 => "0101110011010010", 6982 => "1111101101010011", 6983 => "1011011000011110", 6984 => "0111101001001101", 6985 => "0100110110111000", 6986 => "0001111111011101", 6987 => "1110001011111011", 6988 => "1011000110000101", 6989 => "1010111110011110", 6990 => "1100110110001001", 6991 => "0011101111000111", 6992 => "0010010000111100", 6993 => "0101001110101110", 6994 => "0101110111011111", 6995 => "1000011001001100", 6996 => "0000000001010111", 6997 => "1111000111010100", 6998 => "1110111110110010", 6999 => "0010111111001001", 7000 => "1001100100000100", 7001 => "0011100100010110", 7002 => "0110011001100000", 7003 => "0100110010111111", 7004 => "1111010111110101", 7005 => "1000111001000100", 7006 => "0001110011111100", 7007 => "1101000100011010", 7008 => "0011010101011001", 7009 => "0101111000011010", 7010 => "1000000110101011", 7011 => "0101000011101001", 7012 => "1111101111011110", 7013 => "1111011111011110", 7014 => "1010110001110011", 7015 => "0010000100000110", 7016 => "1000100010110110", 7017 => "0000110101010100", 7018 => "0011001100001010", 7019 => "0101100111000001", 7020 => "0111100100010100", 7021 => "1100010000001100", 7022 => "0101010000110110", 7023 => "0101011011000011", 7024 => "1000111011101010", 7025 => "0111101110001001", 7026 => "1011000001111111", 7027 => "1011111101001011", 7028 => "1101000100110111", 7029 => "1011110010011011", 7030 => "1010010001001000", 7031 => "0010111111011000", 7032 => "0111100000010100", 7033 => "0110111100111100", 7034 => "0100001111100110", 7035 => "0101101001111010", 7036 => "0001111010101111", 7037 => "1100101100010110", 7038 => "1000011011110110", 7039 => "0110011010001110", 7040 => "1000111110000111", 7041 => "0011011100000101", 7042 => "1010001110010101", 7043 => "1100000110100111", 7044 => "0011000010000011", 7045 => "1101101000110110", 7046 => "1101101001101111", 7047 => "1001101110110010", 7048 => "0101001101000101", 7049 => "0101000111001110", 7050 => "0010010010000011", 7051 => "0100011100010111", 7052 => "0101100001001011", 7053 => "1110000010010100", 7054 => "0010001111000111", 7055 => "0000011001011011", 7056 => "1000001101100100", 7057 => "0010000110100000", 7058 => "0000000011101111", 7059 => "1000101011111111", 7060 => "0010100100100011", 7061 => "0110000110000110", 7062 => "0110000101011100", 7063 => "0001110101000001", 7064 => "0000010100001010", 7065 => "1101001101001100", 7066 => "0101010101010101", 7067 => "1110111010110110", 7068 => "0100000100000100", 7069 => "0001000001000111", 7070 => "1110111101110010", 7071 => "1001101011100000", 7072 => "0000000000011011", 7073 => "1110100110100111", 7074 => "0110101100110010", 7075 => "1111001101010000", 7076 => "0111011010001111", 7077 => "1000001111111000", 7078 => "1000001010100000", 7079 => "0011111000000010", 7080 => "1001000100010100", 7081 => "1111100101011100", 7082 => "1000100100101100", 7083 => "0100100001010010", 7084 => "1110111111101011", 7085 => "0010111011100000", 7086 => "0011110010011011", 7087 => "0010000111101111", 7088 => "1010110111001000", 7089 => "1111101101011100", 7090 => "0001010110100000", 7091 => "0101000100101001", 7092 => "1100011100100001", 7093 => "1100000011100100", 7094 => "0110111010110011", 7095 => "1011001010000001", 7096 => "0000101101011110", 7097 => "0001000111011000", 7098 => "1001010011100101", 7099 => "0001010011100101", 7100 => "0001001100110011", 7101 => "1101101101011000", 7102 => "1110100011100000", 7103 => "1100101110111011", 7104 => "1000000110111010", 7105 => "1001000000001100", 7106 => "1111100000101101", 7107 => "0100001011110001", 7108 => "0010001001101111", 7109 => "1101010000101011", 7110 => "0000100010011000", 7111 => "0101111111001100", 7112 => "1101000100001101", 7113 => "0010111110010100", 7114 => "0011100011101100", 7115 => "1011110100110001", 7116 => "0111101100101100", 7117 => "1101111110110111", 7118 => "0000001101101001", 7119 => "1100010101110100", 7120 => "0001101001010101", 7121 => "0111011011110001", 7122 => "1111110000011101", 7123 => "0101000001010110", 7124 => "1001110011100000", 7125 => "0101111100101011", 7126 => "1101000011010110", 7127 => "0100001111110111", 7128 => "1101011101011111", 7129 => "0010010000000010", 7130 => "0011110101100000", 7131 => "0111001110010100", 7132 => "0011000110111100", 7133 => "0000000000011011", 7134 => "0100010101111110", 7135 => "0110111001011101", 7136 => "1110100100010101", 7137 => "0111011000110001", 7138 => "1011011011010010", 7139 => "1010101110001111", 7140 => "1100111000010110", 7141 => "1111100000010001", 7142 => "1101101100001000", 7143 => "0100110010000100", 7144 => "1111000100001110", 7145 => "1010111111101101", 7146 => "0110000001000001", 7147 => "0110110001000101", 7148 => "1101101110000110", 7149 => "1000010101000001", 7150 => "0010101010111110", 7151 => "0000010000101100", 7152 => "1110100001010001", 7153 => "1101100010010000", 7154 => "0011010100011011", 7155 => "1001110111111111", 7156 => "1000010110100100", 7157 => "1011000001011010", 7158 => "0111101001010010", 7159 => "1010110110010010", 7160 => "0001001010010111", 7161 => "1111000001101110", 7162 => "1101100101101001", 7163 => "0001000110001000", 7164 => "0010111111100101", 7165 => "1110011011001101", 7166 => "0111110110011101", 7167 => "0111001011010001", 7168 => "1101100111000011", 7169 => "1101010110110110", 7170 => "1000001100101000", 7171 => "0110010000101000", 7172 => "0000100010111111", 7173 => "0010001110100000", 7174 => "0110101000011001", 7175 => "1010110001100001", 7176 => "0101010011110101", 7177 => "0010101000110101", 7178 => "1101011000101011", 7179 => "0111000010011101", 7180 => "0010100101101110", 7181 => "1111001100000110", 7182 => "1110001100111011", 7183 => "1101011010111000", 7184 => "0010110100000110", 7185 => "1011100001100001", 7186 => "0101001111010100", 7187 => "0111110100001100", 7188 => "1110000011110001", 7189 => "1000010011011100", 7190 => "1101010101000111", 7191 => "1010011000011000", 7192 => "0111000100001100", 7193 => "0100111001100011", 7194 => "1101110011100101", 7195 => "0000110011010011", 7196 => "1100111010100001", 7197 => "0010111010100101", 7198 => "1001100100010010", 7199 => "1101010001100000", 7200 => "0100010100000100", 7201 => "0100101000001000", 7202 => "0010101101101110", 7203 => "1101101011100010", 7204 => "0100100100000011", 7205 => "0101011110000010", 7206 => "0101101010110001", 7207 => "1011010001011001", 7208 => "0111110010001110", 7209 => "0111000011100101", 7210 => "0100000011110111", 7211 => "0100111100011100", 7212 => "0110101011101000", 7213 => "1100011101100111", 7214 => "1001010110001100", 7215 => "1010011001111011", 7216 => "1110011111010110", 7217 => "0001111011111001", 7218 => "0100110101101101", 7219 => "0111101111111110", 7220 => "0100001001100001", 7221 => "1110000010011111", 7222 => "1001101010001100", 7223 => "1000111001111101", 7224 => "0001111110110011", 7225 => "1011010100101001", 7226 => "0111011000100100", 7227 => "0011001100100001", 7228 => "0001001010011111", 7229 => "0010010001111110", 7230 => "0100011100010110", 7231 => "0010011101001100", 7232 => "0000011000100101", 7233 => "0100101001100000", 7234 => "1110000010101011", 7235 => "0000110010110001", 7236 => "1010011111100110", 7237 => "0100000001110010", 7238 => "1111101010111011", 7239 => "1110000101010110", 7240 => "0100111100110001", 7241 => "0111011001101011", 7242 => "0110010111011100", 7243 => "0010001011010011", 7244 => "0000000000110000", 7245 => "1110100001001010", 7246 => "1111110010111111", 7247 => "1111011110111101", 7248 => "0100011101101010", 7249 => "1000011100101110", 7250 => "0111011000010101", 7251 => "0111100011111001", 7252 => "0010111001111100", 7253 => "0001100011001101", 7254 => "1010101000001101", 7255 => "1011001000100101", 7256 => "1111010011001110", 7257 => "1010100100110000", 7258 => "0011100110000010", 7259 => "0100101010011010", 7260 => "0000000010001011", 7261 => "0011101100000010", 7262 => "0100110011101110", 7263 => "1000111011010000", 7264 => "0100001001001101", 7265 => "0101110111010010", 7266 => "1011011110000000", 7267 => "1000011111010010", 7268 => "0101100111000001", 7269 => "1110010110101110", 7270 => "1101111101011000", 7271 => "0101000100111000", 7272 => "1011000101100001", 7273 => "0100000101000001", 7274 => "1110001101111001", 7275 => "1111111101100110", 7276 => "1111100111110001", 7277 => "0010111001110001", 7278 => "1000101101010010", 7279 => "1011111010101101", 7280 => "0001100100101010", 7281 => "1010101000100101", 7282 => "0100100000100000", 7283 => "0100011110110101", 7284 => "1100101010010101", 7285 => "1100000100111000", 7286 => "1001110000101001", 7287 => "1100010111100000", 7288 => "0111111001010011", 7289 => "1010010111000101", 7290 => "0101100101111110", 7291 => "1100000100001000", 7292 => "1001011110110110", 7293 => "0101110000011010", 7294 => "1101001111101011", 7295 => "1111111110000001", 7296 => "0100111011101110", 7297 => "0001111111000001", 7298 => "1110101010101010", 7299 => "1110010011001100", 7300 => "1000101100000000", 7301 => "0001111000110001", 7302 => "0100110100111111", 7303 => "1101100001010010", 7304 => "0101111111100111", 7305 => "0011001110100111", 7306 => "1101111010100010", 7307 => "0101101101101111", 7308 => "1011000110001101", 7309 => "1100001101011000", 7310 => "1000110000001000", 7311 => "0101100011010110", 7312 => "1111111111010100", 7313 => "1101011100111011", 7314 => "0101101000110011", 7315 => "0101101110111010", 7316 => "0001111111111101", 7317 => "0111100001110100", 7318 => "0010110011001011", 7319 => "1001101011110111", 7320 => "1010001011101111", 7321 => "0010011011000101", 7322 => "1001110101110100", 7323 => "1111110111111110", 7324 => "0111001000100010", 7325 => "0001110000001101", 7326 => "0010111010000010", 7327 => "1111101110001110", 7328 => "1010010111001011", 7329 => "0010001011010100", 7330 => "1101001010011000", 7331 => "1101110010110001", 7332 => "1101110001100001", 7333 => "1100101010010000", 7334 => "0110010110110101", 7335 => "0000110100100111", 7336 => "0111011001001011", 7337 => "1000110110101010", 7338 => "1100010111110010", 7339 => "1100100000000000", 7340 => "1000101010111011", 7341 => "1000011000001100", 7342 => "0000111010110000", 7343 => "1110100101010000", 7344 => "1001101000011011", 7345 => "0111010010010010", 7346 => "0110111000000110", 7347 => "1010011100000010", 7348 => "1101001111111110", 7349 => "1001110010100110", 7350 => "0010101101011001", 7351 => "0011101001111011", 7352 => "1000010000100101", 7353 => "1110000111100001", 7354 => "1001101001101010", 7355 => "1101100000111010", 7356 => "0111010101100010", 7357 => "1100101101001101", 7358 => "1001100110101000", 7359 => "1110101011101011", 7360 => "1101101101000101", 7361 => "1001000101000101", 7362 => "0100111100100101", 7363 => "1101111100110101", 7364 => "1000000110000000", 7365 => "0000010111101001", 7366 => "1010000000011001", 7367 => "0111111101000100", 7368 => "1110000101011101", 7369 => "1101110011001110", 7370 => "0100011001111101", 7371 => "1111010011010111", 7372 => "1101001101101110", 7373 => "1111111010000010", 7374 => "0001110010000001", 7375 => "0111110111101011", 7376 => "1100011001010111", 7377 => "0000011010100010", 7378 => "1110101100011111", 7379 => "0000010100101100", 7380 => "0100111000011001", 7381 => "0111000010001010", 7382 => "1101011101101101", 7383 => "0111111001001010", 7384 => "0000011011001111", 7385 => "0001000001001000", 7386 => "1100110010010000", 7387 => "0101001010011010", 7388 => "1010001011101111", 7389 => "1011010001000001", 7390 => "0111111011100000", 7391 => "1101011110110000", 7392 => "0010000000100011", 7393 => "0101010001110010", 7394 => "1100101100100001", 7395 => "0000111101111001", 7396 => "0100111001010011", 7397 => "1000000011111010", 7398 => "0001010000101010", 7399 => "1101110001100000", 7400 => "0100001000110011", 7401 => "0011000000010100", 7402 => "1011100111001101", 7403 => "0010111110111110", 7404 => "1111011101100101", 7405 => "0000001000110101", 7406 => "1010011101000000", 7407 => "1101000111011011", 7408 => "1000000110010101", 7409 => "1100011111000101", 7410 => "1010100001111111", 7411 => "0010110011001001", 7412 => "1101011011101100", 7413 => "0101101010101101", 7414 => "0000010110110010", 7415 => "1000001101101000", 7416 => "1011001110110011", 7417 => "1000110110100111", 7418 => "1111011111101110", 7419 => "1100011101100010", 7420 => "1110100010000000", 7421 => "0101111100101010", 7422 => "1000011101111001", 7423 => "0011010100000011", 7424 => "0011000010011111", 7425 => "0001110001000001", 7426 => "1010000000000110", 7427 => "1101110010100111", 7428 => "1010010101111011", 7429 => "1101001100001000", 7430 => "1011011000000000", 7431 => "1000001101000000", 7432 => "1101000110010001", 7433 => "0000001101100010", 7434 => "1000011111101001", 7435 => "0100101110111010", 7436 => "0100110001001001", 7437 => "1110110011011111", 7438 => "1010011101101010", 7439 => "0101000110010011", 7440 => "0010101010000100", 7441 => "1100011000101100", 7442 => "0011001110011100", 7443 => "0010010100011101", 7444 => "1010100000110100", 7445 => "1000000110110010", 7446 => "0111101111101111", 7447 => "0000101011000001", 7448 => "1111100111110101", 7449 => "0101011011100100", 7450 => "0000000100001010", 7451 => "1010011001100101", 7452 => "0110100110101101", 7453 => "1000101110001100", 7454 => "1101010010101001", 7455 => "1000101000000110", 7456 => "0101100000101111", 7457 => "1110110010001001", 7458 => "0000101100100110", 7459 => "0010110110011010", 7460 => "1001100110000011", 7461 => "1100100110010101", 7462 => "1001111010000101", 7463 => "0101011111101100", 7464 => "0000001010111111", 7465 => "1111111000100101", 7466 => "0000001010100110", 7467 => "1000011011111000", 7468 => "0100101000000111", 7469 => "1110101001110110", 7470 => "0110011011000111", 7471 => "0110100010011100", 7472 => "1011001010000111", 7473 => "1101100110011010", 7474 => "0100011011111110", 7475 => "0011001011001011", 7476 => "1111011110011001", 7477 => "1011100011100111", 7478 => "1110100111100101", 7479 => "1001101000010101", 7480 => "1011101110001100", 7481 => "1011101111110001", 7482 => "1111110101110000", 7483 => "0111101001001111", 7484 => "0000001000011101", 7485 => "1010011110001100", 7486 => "0000111110101011", 7487 => "1000111010011100", 7488 => "1101111110010111", 7489 => "1011010110001101", 7490 => "1100111110010011", 7491 => "0110100001010111", 7492 => "1011001000101011", 7493 => "0000110100001111", 7494 => "1011000001000000", 7495 => "1011101010100001", 7496 => "1111010001011111", 7497 => "0011100100010111", 7498 => "1110111001111010", 7499 => "1110110011100011", 7500 => "1111010000000001", 7501 => "0110001000011101", 7502 => "1010110100101100", 7503 => "0010101100101000", 7504 => "0100111100100010", 7505 => "0011111100101000", 7506 => "0000001011001111", 7507 => "1111101011010110", 7508 => "0001101000010110", 7509 => "0100000000001001", 7510 => "0100011101101011", 7511 => "1010001011100001", 7512 => "0001010110010111", 7513 => "1110010010101011", 7514 => "0010110001101001", 7515 => "0110010101010010", 7516 => "0011011010100111", 7517 => "0011100011100010", 7518 => "1000011100010010", 7519 => "1101111001111001", 7520 => "1100010101100010", 7521 => "1101110100100010", 7522 => "1100100111100010", 7523 => "0110010000000110", 7524 => "1100011001010010", 7525 => "0011110110110111", 7526 => "0000001111000011", 7527 => "1100101111010010", 7528 => "1010010100000100", 7529 => "1001010010100110", 7530 => "0110001001101011", 7531 => "0001001010100110", 7532 => "1110010000101011", 7533 => "0000000010011111", 7534 => "0010111110110110", 7535 => "0001000100100110", 7536 => "1001001010001101", 7537 => "0000110010100000", 7538 => "1000100011011000", 7539 => "1111111010011101", 7540 => "1100111111011111", 7541 => "0100111010011000", 7542 => "1111010011000001", 7543 => "1010110011000000", 7544 => "0111101001011000", 7545 => "0101011000010001", 7546 => "0100100001111000", 7547 => "0001001001001000", 7548 => "0101000011111001", 7549 => "1110110000110111", 7550 => "0010110110001011", 7551 => "1010100111011110", 7552 => "0000011111010101", 7553 => "1100001001010010", 7554 => "1010110101010100", 7555 => "0010000100110100", 7556 => "1011110100100000", 7557 => "0111000001001100", 7558 => "1100001111001100", 7559 => "0111010010100111", 7560 => "0100001101000100", 7561 => "0010011001100011", 7562 => "1010001110101000", 7563 => "0010010101100000", 7564 => "0010111000111100", 7565 => "0111110000001111", 7566 => "0000110000100110", 7567 => "1101100101000100", 7568 => "1110101010011110", 7569 => "0111001100001000", 7570 => "1110100000000000", 7571 => "1100101111000010", 7572 => "0100111010000001", 7573 => "0010111111011101", 7574 => "1001100001000001", 7575 => "1010111011011010", 7576 => "1011011100110001", 7577 => "0111010111111000", 7578 => "0101100001111010", 7579 => "1111110101001110", 7580 => "1011011011111001", 7581 => "0111101100010010", 7582 => "0000011001111010", 7583 => "1011010101111111", 7584 => "0101110001000111", 7585 => "0001101101100111", 7586 => "1101100111111011", 7587 => "1001100111000100", 7588 => "1101011010101100", 7589 => "0001001010100010", 7590 => "0011011110101011", 7591 => "0100000001111010", 7592 => "1010110001000011", 7593 => "0001101100101001", 7594 => "0000110001101101", 7595 => "1010110111001010", 7596 => "0101100011000101", 7597 => "0100010010000010", 7598 => "0111000101111111", 7599 => "0011111101110101", 7600 => "0010111110000100", 7601 => "0001101111000100", 7602 => "1000001001010100", 7603 => "0110111101011100", 7604 => "0101111111110110", 7605 => "0101101001101001", 7606 => "1100100000110011", 7607 => "0111010110101000", 7608 => "1110110001100011", 7609 => "0101110100110111", 7610 => "1011001111001011", 7611 => "0100001011000000", 7612 => "1001001011010111", 7613 => "0101001111011010", 7614 => "0110000110101010", 7615 => "1011010111100110", 7616 => "1011101111011100", 7617 => "1110101111001101", 7618 => "1100001101000010", 7619 => "0100010011000000", 7620 => "0100111000010001", 7621 => "1000000001110111", 7622 => "1000111010101110", 7623 => "1010000001001001", 7624 => "1010010000100011", 7625 => "1010000001100110", 7626 => "0110001001101110", 7627 => "0110100010001111", 7628 => "1000001010101111", 7629 => "0100001010000100", 7630 => "1110000000010000", 7631 => "0111101000011000", 7632 => "0101100111010011", 7633 => "1011110101100111", 7634 => "0011000100010100", 7635 => "0000001111101000", 7636 => "1001111011010011", 7637 => "0011100110110101", 7638 => "0111000011111001", 7639 => "0100010001011110", 7640 => "0110110000100101", 7641 => "1111000011001110", 7642 => "0101110111001011", 7643 => "1110101101011100", 7644 => "1001010100110111", 7645 => "1010101010110001", 7646 => "1100101111000000", 7647 => "1110111010101110", 7648 => "1101101101101011", 7649 => "0110011100000110", 7650 => "1100111100100001", 7651 => "1000101010010010", 7652 => "0110110111110000", 7653 => "1000011100100000", 7654 => "0111001000010101", 7655 => "1110001000101011", 7656 => "0111011011010011", 7657 => "0011101011010100", 7658 => "0011010101100101", 7659 => "0010011011101000", 7660 => "1010000100111010", 7661 => "0010000111100110", 7662 => "0000110011111101", 7663 => "1101010110010001", 7664 => "0001011010010110", 7665 => "1010100011101111", 7666 => "1010101001000010", 7667 => "0010100101110100", 7668 => "1100001111111101", 7669 => "0010001101001110", 7670 => "0010011100111110", 7671 => "1011001010000111", 7672 => "1100010001001001", 7673 => "1101000000011011", 7674 => "1101110001111000", 7675 => "0001010011001101", 7676 => "1010110100100011", 7677 => "0001101011000101", 7678 => "1100010100110100", 7679 => "0011000101011001", 7680 => "1101100011101001", 7681 => "1111101101100110", 7682 => "1010110110011110", 7683 => "1110001111000111", 7684 => "1010101001010100", 7685 => "0011011111110011", 7686 => "0011101100110110", 7687 => "1100111100000011", 7688 => "1101100000011101", 7689 => "1110010011000001", 7690 => "1011101000110001", 7691 => "0110010111100111", 7692 => "1100011100111000", 7693 => "0011011010111001", 7694 => "1100100100000011", 7695 => "1001110100000010", 7696 => "0000101011100110", 7697 => "1001010111100110", 7698 => "0100010100001111", 7699 => "1111011010100101", 7700 => "0100001100100000", 7701 => "1011101010000100", 7702 => "1110111111011111", 7703 => "1000101101001000", 7704 => "0010110010101010", 7705 => "0110101001001001", 7706 => "1101010110011111", 7707 => "0001100101011001", 7708 => "1010100101001001", 7709 => "0111010111101110", 7710 => "0101010000001000", 7711 => "0011100011111110", 7712 => "1001111111110001", 7713 => "0101011000101100", 7714 => "1011111000110101", 7715 => "1101101000001110", 7716 => "0010011011000001", 7717 => "1101101011111011", 7718 => "1011100000001001", 7719 => "1001101101011110", 7720 => "1110000010000110", 7721 => "0111110011001000", 7722 => "0011110011011101", 7723 => "0101000100000001", 7724 => "1101011011111111", 7725 => "1101110010111100", 7726 => "0010101000011101", 7727 => "1000101011010101", 7728 => "1111011010110111", 7729 => "1010110110010100", 7730 => "0101000101100110", 7731 => "1011000010100100", 7732 => "1100001010011111", 7733 => "1010101110110111", 7734 => "0101111000110010", 7735 => "1101101011010111", 7736 => "1100101011001100", 7737 => "1001111000111100", 7738 => "0110110001000001", 7739 => "0011101010001100", 7740 => "0110011100000000", 7741 => "0110110110001000", 7742 => "1110011000100001", 7743 => "0100111000111000", 7744 => "1101011100011010", 7745 => "0000000110101110", 7746 => "0000111000000100", 7747 => "0111100111111001", 7748 => "1010000111100010", 7749 => "0010100110001001", 7750 => "1011011001011011", 7751 => "0010011011000110", 7752 => "1111101100001010", 7753 => "0100011001111110", 7754 => "1001011100000010", 7755 => "1000010101100010", 7756 => "1001011011101011", 7757 => "1011111101111110", 7758 => "0001010000100010", 7759 => "1000111110101101", 7760 => "1100010010100100", 7761 => "0000111111011010", 7762 => "1100001101110111", 7763 => "0000001010011001", 7764 => "1010001000100100", 7765 => "0010110111000111", 7766 => "0010101000001100", 7767 => "1000101001111111", 7768 => "1110010110000101", 7769 => "0100101000101000", 7770 => "1100010010011001", 7771 => "0100011010000011", 7772 => "1101011010110000", 7773 => "0110011111110010", 7774 => "0110000001011001", 7775 => "0110101110101101", 7776 => "1011011000101010", 7777 => "1010001011001010", 7778 => "1110011111000101", 7779 => "1010010110011010", 7780 => "1011111010010110", 7781 => "1001110100001100", 7782 => "0101001111001000", 7783 => "1101111111011010", 7784 => "1110011100010001", 7785 => "0001011111100100", 7786 => "0100001100010100", 7787 => "0000111010001001", 7788 => "1111000011101001", 7789 => "1111011011010110", 7790 => "1111011001111000", 7791 => "0011011110101110", 7792 => "0100110110000011", 7793 => "0010011011110000", 7794 => "1100000010101001", 7795 => "0101111111100001", 7796 => "0011111010110000", 7797 => "0000010001001000", 7798 => "0100000110000111", 7799 => "0000000000100000", 7800 => "1001001010001110", 7801 => "0001000000100100", 7802 => "1111110000110100", 7803 => "1000110110101111", 7804 => "1111100111001001", 7805 => "1011100010001110", 7806 => "0010100111101100", 7807 => "0000111010101101", 7808 => "0010110101010010", 7809 => "1111100010000001", 7810 => "0001010111010011", 7811 => "0100111100001011", 7812 => "0001100100010001", 7813 => "1100110100101110", 7814 => "1011000010111111", 7815 => "0000110111110010", 7816 => "1110101000011111", 7817 => "0010000011001010", 7818 => "1100101011010001", 7819 => "1011110000000000", 7820 => "1101000101101000", 7821 => "0011101110001111", 7822 => "1001001111101011", 7823 => "1001001111100001", 7824 => "0101110100110011", 7825 => "0011111010110010", 7826 => "0100111011001010", 7827 => "0000010000001001", 7828 => "1011100001011011", 7829 => "0001001000011000", 7830 => "0000110011100110", 7831 => "1110100000000011", 7832 => "0010111111100011", 7833 => "0000110011010100", 7834 => "1110001111101000", 7835 => "1001011100111011", 7836 => "0001101101100011", 7837 => "0011010001100011", 7838 => "1100101001111000", 7839 => "1000100101011010", 7840 => "1011001010110100", 7841 => "1110010110110110", 7842 => "1110111010001101", 7843 => "0110101100101101", 7844 => "1110100101011111", 7845 => "0011110010111110", 7846 => "1011111110000110", 7847 => "1001000011010100", 7848 => "0001001111011001", 7849 => "1110100111010100", 7850 => "1001010011111010", 7851 => "0011001011111001", 7852 => "0000110011111001", 7853 => "1010001010000011", 7854 => "1010101010100110", 7855 => "1100111010111000", 7856 => "0110111001010101", 7857 => "0100000010000010", 7858 => "1101100100001001", 7859 => "0101000011111110", 7860 => "0100100011110010", 7861 => "1110100110110101", 7862 => "0010010111011000", 7863 => "1100011110001101", 7864 => "1011100001101101", 7865 => "1100100011000100", 7866 => "1111110001001010", 7867 => "1001111011100010", 7868 => "0011111100100110", 7869 => "1000011101100010", 7870 => "0011110101000000", 7871 => "0100101010110000", 7872 => "0100111010110001", 7873 => "1101011010111010", 7874 => "0111001101000100", 7875 => "1111000110001101", 7876 => "0110011101101001", 7877 => "1100010100111101", 7878 => "1000011010011001", 7879 => "0111001000111011", 7880 => "1101101101110001", 7881 => "1000111010111101", 7882 => "0001111001101100", 7883 => "1011101110010110", 7884 => "0010100000110011", 7885 => "1010011101001001", 7886 => "1001100011001101", 7887 => "1110111110101101", 7888 => "1110001100100001", 7889 => "0100001001000010", 7890 => "0101100011000010", 7891 => "1110001010101001", 7892 => "0010100110000001", 7893 => "0110011000000011", 7894 => "1101101001000001", 7895 => "0100100101110000", 7896 => "0001111010011100", 7897 => "1110001101100110", 7898 => "1110100101010010", 7899 => "0111000110000011", 7900 => "1010000110010011", 7901 => "1001111001110011", 7902 => "1011101011101101", 7903 => "0110100111011101", 7904 => "1110110100110100", 7905 => "0011000010001110", 7906 => "0000101011011110", 7907 => "1001010001110111", 7908 => "0011011110010100", 7909 => "1001010000000010", 7910 => "0111011111010000", 7911 => "1011100010111010", 7912 => "1110000110011000", 7913 => "0111011101010111", 7914 => "1100000110011110", 7915 => "1110010010011111", 7916 => "0100110011011010", 7917 => "0101101101011011", 7918 => "0000111000011101", 7919 => "1100100000000100", 7920 => "0110101000101101", 7921 => "1011011001001001", 7922 => "1110001110001100", 7923 => "1010001001111000", 7924 => "0011011010001001", 7925 => "1100100101011101", 7926 => "0101100010000010", 7927 => "0001000011111110", 7928 => "1100001101100111", 7929 => "0100110010000101", 7930 => "0011111001101000", 7931 => "1000001001100011", 7932 => "1110010111110101", 7933 => "0101100001010010", 7934 => "0111100011010011", 7935 => "1011001100000111", 7936 => "0001001000110001", 7937 => "0111110101101100", 7938 => "0100011010001101", 7939 => "0000000011110100", 7940 => "1000001010101011", 7941 => "1011001011011001", 7942 => "1000000011100111", 7943 => "0111101111010001", 7944 => "1101001001101110", 7945 => "1111011101110101", 7946 => "0011001001100000", 7947 => "0100000111000111", 7948 => "1110101111110111", 7949 => "0001000010000100", 7950 => "0000001001100110", 7951 => "0010000100110101", 7952 => "0110010111010000", 7953 => "1111011110100100", 7954 => "1111001011101001", 7955 => "1000001101010100", 7956 => "1111100011111101", 7957 => "0101100001000101", 7958 => "0011101000001011", 7959 => "0110010000100110", 7960 => "0010001000101001", 7961 => "1101001000010011", 7962 => "1110001000111000", 7963 => "1000110111010011", 7964 => "1000111000011111", 7965 => "0111101100101111", 7966 => "0000100110011110", 7967 => "1110001101100110", 7968 => "1001001000011011", 7969 => "0111001111011010", 7970 => "1011001101000010", 7971 => "1010000001100100", 7972 => "0001001101100011", 7973 => "0000001111010100", 7974 => "1011100111111000", 7975 => "1011001001010110", 7976 => "0101010000010101", 7977 => "0111101101101011", 7978 => "1010010110010110", 7979 => "0010100000000111", 7980 => "0101110110010000", 7981 => "0001100110110010", 7982 => "0100010010001111", 7983 => "0100100011011001", 7984 => "0111101001111111", 7985 => "0000110100111111", 7986 => "1111000011101110", 7987 => "1011001010010011", 7988 => "1001110000101001", 7989 => "0100010110010111", 7990 => "1110010100010110", 7991 => "0011000000100111", 7992 => "1111110011110101", 7993 => "0010010110110100", 7994 => "0111011010011010", 7995 => "0010101011001010", 7996 => "0000110100111001", 7997 => "0110101010001111", 7998 => "1110101110000110", 7999 => "1111000100000101", 8000 => "0010110101110101", 8001 => "0111101011100011", 8002 => "0000110000011000", 8003 => "0001001000100000", 8004 => "1001010001000011", 8005 => "1011101111011111", 8006 => "0010110011001010", 8007 => "0011000001101111", 8008 => "1011010001110100", 8009 => "0011111101000011", 8010 => "1001100011110011", 8011 => "1101010001110111", 8012 => "0101000111011000", 8013 => "1011000111001001", 8014 => "1001111101000010", 8015 => "0000010100111101", 8016 => "1100110100001111", 8017 => "0110010101101111", 8018 => "1010010110100001", 8019 => "0000010110001101", 8020 => "0000001111001000", 8021 => "0100011001011001", 8022 => "0111001100001001", 8023 => "1100000111010100", 8024 => "1000000000100111", 8025 => "0100101010100001", 8026 => "1111011000001010", 8027 => "0011100100011100", 8028 => "1010111001110111", 8029 => "1110011011100111", 8030 => "1000100010001000", 8031 => "0011000111001011", 8032 => "0101101100110010", 8033 => "1101001110100101", 8034 => "1001100111101010", 8035 => "1110001000101111", 8036 => "0100001101111001", 8037 => "0111100111110010", 8038 => "0110100011001001", 8039 => "0100001011010111", 8040 => "0111110110111001", 8041 => "1000110110011100", 8042 => "0001011000100001", 8043 => "0110101101010010", 8044 => "0010101100110101", 8045 => "1110111101111001", 8046 => "0101111010000101", 8047 => "0101101011011100", 8048 => "0111110110110011", 8049 => "0000011001110101", 8050 => "0010011111011111", 8051 => "0000101010000001", 8052 => "0000100011100110", 8053 => "1000011110101001", 8054 => "1000011101011000", 8055 => "0010101010100000", 8056 => "1101000110010101", 8057 => "0101110100000011", 8058 => "1010110101111110", 8059 => "0001101011101010", 8060 => "1010011111001101", 8061 => "1110000110110011", 8062 => "0110011000001010", 8063 => "1011011100010001", 8064 => "0111001000110111", 8065 => "0010011110110111", 8066 => "0110000110000000", 8067 => "1010111000000000", 8068 => "1001001101111111", 8069 => "1000100100111000", 8070 => "1111100000011111", 8071 => "1000000001110100", 8072 => "0000101000010001", 8073 => "0101010110001100", 8074 => "0010110010000101", 8075 => "1111101000100110", 8076 => "0111011001011001", 8077 => "1110001101101101", 8078 => "0101100000001000", 8079 => "0101000101010010", 8080 => "1001010101001110", 8081 => "1001110100110100", 8082 => "1010001010101001", 8083 => "1100000110100001", 8084 => "1010001101000100", 8085 => "0100101001100110", 8086 => "1000111110111011", 8087 => "0010100101110000", 8088 => "1110110101111111", 8089 => "0000011000101100", 8090 => "1111101110000101", 8091 => "0001000000101001", 8092 => "1001110010101101", 8093 => "0110100010010100", 8094 => "1010111011111100", 8095 => "0000110111110001", 8096 => "0111001111010111", 8097 => "1100111010100100", 8098 => "1000000110000001", 8099 => "0101011101110111", 8100 => "1011011011001001", 8101 => "0111010111000100", 8102 => "1100101100100100", 8103 => "0001010001000111", 8104 => "0110100011101011", 8105 => "1101111100001101", 8106 => "1110101000100010", 8107 => "0010111011101100", 8108 => "1111100111111111", 8109 => "1101000000010000", 8110 => "0001101111100011", 8111 => "1001000101011100", 8112 => "0110010110010010", 8113 => "1010011011001100", 8114 => "0000010111001001", 8115 => "1001000101101001", 8116 => "1110000101011000", 8117 => "0110110000111100", 8118 => "0011001001110100", 8119 => "1100110001101111", 8120 => "1101100011000101", 8121 => "0000001101001110", 8122 => "1110101001101100", 8123 => "0000000100001100", 8124 => "1110001000111100", 8125 => "1000101101100010", 8126 => "1000110110001101", 8127 => "0000011100111000", 8128 => "1110001010101001", 8129 => "0110000010111001", 8130 => "0010111111100110", 8131 => "1110100001001000", 8132 => "1011000011011001", 8133 => "0000111010011010", 8134 => "0110101101000110", 8135 => "1110111001111101", 8136 => "1111011110000100", 8137 => "1111001101010111", 8138 => "1000011011010100", 8139 => "1101000001010100", 8140 => "1111010001110111", 8141 => "1000101100111010", 8142 => "1101011011111000", 8143 => "0111000100001111", 8144 => "1100100110011010", 8145 => "1011001000100011", 8146 => "0000000111011101", 8147 => "0110110011100001", 8148 => "1001000110000111", 8149 => "0101000101100001", 8150 => "0110111011001111", 8151 => "0101111011000100", 8152 => "0101001110101100", 8153 => "1110100000000110", 8154 => "1010000100001101", 8155 => "1111001100010000", 8156 => "0101010011101101", 8157 => "0000001100000000", 8158 => "1011110110101001", 8159 => "1111111111000001", 8160 => "1101011111011011", 8161 => "0111000111111001", 8162 => "1000001111100100", 8163 => "0110001011011100", 8164 => "1100110000001111", 8165 => "0010001100110010", 8166 => "1000110001001010", 8167 => "0111011001101101", 8168 => "0001101100111111", 8169 => "0001011010101100", 8170 => "0011011111111011", 8171 => "0011011011000100", 8172 => "1001110010001001", 8173 => "1110000111110111", 8174 => "1011001100001001", 8175 => "0000010010111111", 8176 => "0010111011101110", 8177 => "0101000001101110", 8178 => "1110010110111101", 8179 => "0001001001100110", 8180 => "0100111011101010", 8181 => "1110000010101111", 8182 => "1101110101011110", 8183 => "1000011110110100", 8184 => "0101011110111101", 8185 => "1000000100101001", 8186 => "1101111100000111", 8187 => "1110011010101001", 8188 => "1111001001011110", 8189 => "1010101111111010", 8190 => "1111001111010100", 8191 => "1000111010011110", 8192 => "0101100100100010", 8193 => "0001101100100111", 8194 => "0110000000010111", 8195 => "1011100101011010", 8196 => "0001100000111001", 8197 => "0110011111101101", 8198 => "0111000000000011", 8199 => "0111101010110001", 8200 => "0000001001110011", 8201 => "1101000100011101", 8202 => "1100101100010001", 8203 => "1000110010011001", 8204 => "0100101100110001", 8205 => "1100000010100101", 8206 => "0111101111001010", 8207 => "0000101001110101", 8208 => "1001111011110110", 8209 => "1111001010110001", 8210 => "0110001000011010", 8211 => "1000111101101010", 8212 => "1101010011011011", 8213 => "1111010010101101", 8214 => "1100110101011100", 8215 => "0110110110001010", 8216 => "0010011011100010", 8217 => "1001101010100100", 8218 => "0100101111100011", 8219 => "0010011110011110", 8220 => "1111001101011110", 8221 => "1110110101101000", 8222 => "1101001001111111", 8223 => "0100101000010000", 8224 => "1111011111101101", 8225 => "0101111000101011", 8226 => "1010001101101000", 8227 => "0001110011110011", 8228 => "0001100010011000", 8229 => "1110110111001011", 8230 => "0110000001100111", 8231 => "0100010001110011", 8232 => "0010110011010010", 8233 => "1000110100111110", 8234 => "0011010101001100", 8235 => "1101101001110011", 8236 => "1011010010111001", 8237 => "1000011100001011", 8238 => "0010110100001100", 8239 => "0001100110111111", 8240 => "1001101000000011", 8241 => "1101101110101100", 8242 => "0010101010011011", 8243 => "1111100001100110", 8244 => "0000010000010100", 8245 => "1000110111100111", 8246 => "1011001101101000", 8247 => "0001110001111001", 8248 => "0011011001011000", 8249 => "0001101000111110", 8250 => "0010110111000100", 8251 => "0101001011000000", 8252 => "1111100110011110", 8253 => "1111101001001101", 8254 => "1001010110001000", 8255 => "0101011111111101", 8256 => "1010100110000110", 8257 => "0110110101010011", 8258 => "0100111100010111", 8259 => "0001010101111100", 8260 => "1001111000001111", 8261 => "0100111101111010", 8262 => "1001101000110110", 8263 => "1011000011000011", 8264 => "1011111001100001", 8265 => "1100000010001101", 8266 => "1100111000010010", 8267 => "1111000010011101", 8268 => "1001000010001100", 8269 => "1110100011110111", 8270 => "1100110110111000", 8271 => "1011000110001111", 8272 => "1010001011000011", 8273 => "1100100100000100", 8274 => "1010101011000001", 8275 => "1001001011010111", 8276 => "0011110101001110", 8277 => "0011111000011000", 8278 => "1100100110001100", 8279 => "0100100100010100", 8280 => "0100100101100010", 8281 => "0000010101001110", 8282 => "1100010001001011", 8283 => "1111000110101100", 8284 => "0011101011101101", 8285 => "0111001100101100", 8286 => "0011000111101100", 8287 => "1011011011100011", 8288 => "0110100100010011", 8289 => "1010110101011110", 8290 => "0111000101100001", 8291 => "0011011010010101", 8292 => "1111101010101101", 8293 => "1111101100001010", 8294 => "1000101101000010", 8295 => "0000100010001000", 8296 => "1101101001100010", 8297 => "1101110000000001", 8298 => "1000011110101010", 8299 => "0110000000101110", 8300 => "1010000100101110", 8301 => "1000101110110000", 8302 => "0010100001010000", 8303 => "0001110000101001", 8304 => "1010010100001011", 8305 => "0100001011101101", 8306 => "0000001110100101", 8307 => "0101111010001011", 8308 => "1011111001111010", 8309 => "0011100000111011", 8310 => "0001111011100001", 8311 => "0010111001000111", 8312 => "0011111100001001", 8313 => "0010111011111011", 8314 => "1010101100100010", 8315 => "1110011001011110", 8316 => "1000010110111001", 8317 => "1010001000001101", 8318 => "0101010000010011", 8319 => "0111011011101011", 8320 => "1001001011100011", 8321 => "0001111000000011", 8322 => "1100100100111001", 8323 => "0000101101000010", 8324 => "0001010110010001", 8325 => "1000010010000100", 8326 => "0000000100101001", 8327 => "1111111111110010", 8328 => "0000110000001001", 8329 => "0101011111000101", 8330 => "1000111110001011", 8331 => "0100001000100110", 8332 => "1100001001001001", 8333 => "1100100011111011", 8334 => "0011001010001011", 8335 => "0110000000000010", 8336 => "0110000010101011", 8337 => "0111110010111000", 8338 => "1100110000000100", 8339 => "0000000011111100", 8340 => "1011111010000110", 8341 => "0010001001011011", 8342 => "1011110110011000", 8343 => "1000010010110100", 8344 => "0100100101000010", 8345 => "0011111110100010", 8346 => "1001011110111000", 8347 => "0110111111011010", 8348 => "0010000111100000", 8349 => "0111000001101100", 8350 => "1001100101101110", 8351 => "1000111100100101", 8352 => "0101101001110100", 8353 => "0010011000110011", 8354 => "1011111111110101", 8355 => "0011111000010110", 8356 => "1100011000011111", 8357 => "1011001010100000", 8358 => "1010000111010110", 8359 => "1110101010011011", 8360 => "0011111010111000", 8361 => "0011001011101010", 8362 => "0010001011011100", 8363 => "0011010101000001", 8364 => "0000111111111101", 8365 => "1011101011110101", 8366 => "0001110101101101", 8367 => "1111010100001011", 8368 => "1100101011010101", 8369 => "0010010001111001", 8370 => "0001001001101110", 8371 => "1011110011001101", 8372 => "0010010001111100", 8373 => "0110001100110110", 8374 => "1101101100111111", 8375 => "1000110010010111", 8376 => "0010001000010010", 8377 => "1100000100001001", 8378 => "0100010110111100", 8379 => "0110000011110001", 8380 => "0000100010011011", 8381 => "1110001111010011", 8382 => "1011001101000001", 8383 => "0100000100000101", 8384 => "1001011001101001", 8385 => "0101001111001111", 8386 => "0110100101000111", 8387 => "1110000001111100", 8388 => "0111011011101000", 8389 => "0101101001011111", 8390 => "1110010011111000", 8391 => "1000111111001010", 8392 => "1111011010011100", 8393 => "1110000101010110", 8394 => "1000100001001001", 8395 => "0000001010100000", 8396 => "0100010001010110", 8397 => "0101100100100010", 8398 => "1101111110110001", 8399 => "1100111111011110", 8400 => "1111000110000100", 8401 => "1011011001111100", 8402 => "0101111101100101", 8403 => "1001010111100001", 8404 => "1010101110100100", 8405 => "0110100100010001", 8406 => "0010101111000100", 8407 => "1101010100011000", 8408 => "1111111100111100", 8409 => "0000111101000011", 8410 => "0111000110010011", 8411 => "1010111011110100", 8412 => "0011011100111101", 8413 => "1110011110000101", 8414 => "1010100010111101", 8415 => "1110110010111110", 8416 => "0100110100000101", 8417 => "0001100011100101", 8418 => "0111110111110111", 8419 => "0111011000111110", 8420 => "1000001000001111", 8421 => "0010101000100001", 8422 => "0010100111011101", 8423 => "1101111000010100", 8424 => "0000110011101010", 8425 => "0001110011101010", 8426 => "0110000110110001", 8427 => "0100011001000110", 8428 => "1110000001111100", 8429 => "1111110011001110", 8430 => "1100110000011111", 8431 => "0010011101100110", 8432 => "0001101111011000", 8433 => "0011000010100011", 8434 => "0110011011100010", 8435 => "0001011101110001", 8436 => "1101011010011110", 8437 => "0011000000001001", 8438 => "1111101111010101", 8439 => "1110001010111010", 8440 => "1010100000001011", 8441 => "1101010000111010", 8442 => "1000001011011010", 8443 => "0100100000111001", 8444 => "0010000001000101", 8445 => "1010001011101111", 8446 => "1101001011110100", 8447 => "1101100111001011", 8448 => "1001111100101111", 8449 => "1011100000011110", 8450 => "1001000010111111", 8451 => "1001110000101101", 8452 => "0001000101010000", 8453 => "0000100101111100", 8454 => "1011110001001101", 8455 => "1110110111111100", 8456 => "1011011111001001", 8457 => "1011001100010011", 8458 => "1001000111011000", 8459 => "1110010111011000", 8460 => "1000110110011100", 8461 => "0001000001110100", 8462 => "0101110100010101", 8463 => "0010000101000011", 8464 => "0100111110111000", 8465 => "0100111111101011", 8466 => "1011110111100111", 8467 => "0111000111010110", 8468 => "1011010110010100", 8469 => "0101011101101101", 8470 => "1111101100101110", 8471 => "0100110011011011", 8472 => "1111100001101100", 8473 => "1110010100100101", 8474 => "1110101110101100", 8475 => "1101110010010000", 8476 => "0010110010111100", 8477 => "1100110000011000", 8478 => "1100010110000010", 8479 => "1111110001000100", 8480 => "0001110101110000", 8481 => "0011101111101001", 8482 => "1111100101111001", 8483 => "0000011011011001", 8484 => "0101110000110100", 8485 => "0101011000011010", 8486 => "0100011011011010", 8487 => "1101001101001100", 8488 => "1010001011000010", 8489 => "0010101000000010", 8490 => "1001101001001111", 8491 => "1101100010101111", 8492 => "1011010101010110", 8493 => "1010001011111001", 8494 => "1000100111000011", 8495 => "1111101001011001", 8496 => "1010000001010001", 8497 => "1111011000011110", 8498 => "0000011111011100", 8499 => "0001000010110001", 8500 => "0100100001011101", 8501 => "1100000110110111", 8502 => "0101101100111101", 8503 => "1110000111101000", 8504 => "0110001011101010", 8505 => "1110111010001001", 8506 => "1000011001011011", 8507 => "0011001011001111", 8508 => "1100000101110101", 8509 => "0100011010100000", 8510 => "0100010011001010", 8511 => "0110101010101101", 8512 => "1010010110111100", 8513 => "1001110111011100", 8514 => "1010101111100000", 8515 => "0011010101100111", 8516 => "0001010000101101", 8517 => "0101111010111111", 8518 => "0001110010101111", 8519 => "1001001000011101", 8520 => "0000111100000011", 8521 => "1110100000100111", 8522 => "0001110010100010", 8523 => "0000010101111000", 8524 => "1000000110001011", 8525 => "1011010011010110", 8526 => "1010000000011010", 8527 => "0011110100011110", 8528 => "0010111000001010", 8529 => "1111000011001100", 8530 => "0010010001101000", 8531 => "0100101000110100", 8532 => "0101000101001111", 8533 => "0101111011011000", 8534 => "0101100100001000", 8535 => "0011011110011100", 8536 => "0111000100000011", 8537 => "0111011001011111", 8538 => "0101010000001101", 8539 => "0110100100111011", 8540 => "1101011010100101", 8541 => "1100110111101111", 8542 => "1011100101111111", 8543 => "1001000011101010", 8544 => "1001010001010100", 8545 => "0000110011110000", 8546 => "1000100001010110", 8547 => "0111000111110011", 8548 => "0000111010000000", 8549 => "1100100111001010", 8550 => "0010011000100110", 8551 => "0100111101111000", 8552 => "1011111001110000", 8553 => "0110100100000010", 8554 => "1000101000110010", 8555 => "1100010011011110", 8556 => "1110111110010001", 8557 => "1101001001110001", 8558 => "1111011110010111", 8559 => "0001000100101010", 8560 => "0011111110011111", 8561 => "0110001011010010", 8562 => "0101010110010000", 8563 => "0000011101000001", 8564 => "0001111101000011", 8565 => "1010100000100110", 8566 => "1000110101110110", 8567 => "1100001111000000", 8568 => "1110101111100011", 8569 => "1100011110100101", 8570 => "1011100111001011", 8571 => "1110110001000111", 8572 => "1010111101111001", 8573 => "0101000110100000", 8574 => "0001110000000110", 8575 => "0001001110100111", 8576 => "1000011111011100", 8577 => "1101100110111001", 8578 => "0100110000001110", 8579 => "0101111111110101", 8580 => "0011000000001100", 8581 => "0100001111100110", 8582 => "0100101010101100", 8583 => "1101101011010000", 8584 => "1110001110111001", 8585 => "1011010100011001", 8586 => "1001011100010011", 8587 => "0000111101011010", 8588 => "1010011110000101", 8589 => "1000101101111111", 8590 => "0100001100001001", 8591 => "0001101010010111", 8592 => "0011110100000101", 8593 => "1001011111001100", 8594 => "1101110011110000", 8595 => "0101001010110010", 8596 => "1001011010100011", 8597 => "0001110110010001", 8598 => "1000101011010000", 8599 => "1111010110100001", 8600 => "1010101101000101", 8601 => "0010010111111100", 8602 => "1111100111011010", 8603 => "1110001111110111", 8604 => "0000100001010101", 8605 => "1010111000100110", 8606 => "1011110111010111", 8607 => "0000110011111100", 8608 => "1011111100100101", 8609 => "1011100111111001", 8610 => "1111101111101000", 8611 => "1000110010001011", 8612 => "0110010001010100", 8613 => "1110000111110010", 8614 => "0110111011010100", 8615 => "1100110101110001", 8616 => "0011101101011100", 8617 => "0000110111010101", 8618 => "1110010100001010", 8619 => "1001110111101000", 8620 => "1111100000100111", 8621 => "0000111100100010", 8622 => "0100101001100100", 8623 => "1010101101111100", 8624 => "0100011000011100", 8625 => "1001100011110110", 8626 => "0000000010101000", 8627 => "0000011100010001", 8628 => "1111010110101110", 8629 => "1100111100110000", 8630 => "0010111100110101", 8631 => "0011011010000010", 8632 => "0000001010111011", 8633 => "0010000001111100", 8634 => "0011011000110011", 8635 => "0000000000011010", 8636 => "1100110110011110", 8637 => "1110001100011011", 8638 => "0100101000000000", 8639 => "1100011111100110", 8640 => "0111100111101001", 8641 => "1010111001001000", 8642 => "0000001101000001", 8643 => "1000000001000101", 8644 => "1010000000011011", 8645 => "0011011100010000", 8646 => "0000101100101000", 8647 => "1010001000001000", 8648 => "0010000100010010", 8649 => "0101110000110000", 8650 => "0110110110100110", 8651 => "1010100101010000", 8652 => "0001100101101110", 8653 => "1000001101101100", 8654 => "0100100110111010", 8655 => "1011101111111011", 8656 => "0100100101011110", 8657 => "1101101010011111", 8658 => "1010000000000010", 8659 => "1101101011000001", 8660 => "0101100111111011", 8661 => "1001110110010001", 8662 => "0110001101011011", 8663 => "0110100111001100", 8664 => "0111101110010100", 8665 => "0011001111010000", 8666 => "1110000111011001", 8667 => "0000100100001000", 8668 => "0011000010111010", 8669 => "0101011100100111", 8670 => "0100000010111110", 8671 => "0111011001110111", 8672 => "1010000110100010", 8673 => "0111011011010101", 8674 => "1001111110001111", 8675 => "1000100110001001", 8676 => "0011000101010111", 8677 => "0110100000001001", 8678 => "0001001100100111", 8679 => "1110010110110101", 8680 => "1101111000101000", 8681 => "0010101110010001", 8682 => "1111101000101001", 8683 => "1001001011001010", 8684 => "0011010111000010", 8685 => "1000011010111100", 8686 => "0011110110111000", 8687 => "1011000100100000", 8688 => "1000110110001001", 8689 => "1001011010010000", 8690 => "1100011111110100", 8691 => "1010101110101110", 8692 => "0001000100000010", 8693 => "0111010001110011", 8694 => "1010110100111100", 8695 => "1001001001000000", 8696 => "0111100101110101", 8697 => "0111010100110010", 8698 => "0010001011001010", 8699 => "1010010101100110", 8700 => "1111111010011000", 8701 => "1001111000010110", 8702 => "0000100111101011", 8703 => "0000110010000111", 8704 => "1000011101011001", 8705 => "1111000100110100", 8706 => "1000111011010010", 8707 => "1001000011010110", 8708 => "1001001110001011", 8709 => "1110011000010010", 8710 => "0000110010111001", 8711 => "0011000000110011", 8712 => "0011100011000000", 8713 => "0110010101111100", 8714 => "1011110010010101", 8715 => "1101011101001011", 8716 => "0100111010001100", 8717 => "1001011001101011", 8718 => "1111001011010011", 8719 => "1001110100101001", 8720 => "0100000100111000", 8721 => "0000011000001100", 8722 => "1111011110111011", 8723 => "0001111000110111", 8724 => "1111100000101101", 8725 => "1011000101000000", 8726 => "0001110110100110", 8727 => "1110111000111111", 8728 => "1110111011100101", 8729 => "1111011110011101", 8730 => "1011100000001111", 8731 => "1001000011110111", 8732 => "1100011001111001", 8733 => "0000010111001010", 8734 => "0100100001001110", 8735 => "1110100111010111", 8736 => "1010100111010110", 8737 => "0111100010100010", 8738 => "1100001110010111", 8739 => "1100101111111101", 8740 => "0100110110011001", 8741 => "1010001110111001", 8742 => "0010000100110010", 8743 => "0010100001111001", 8744 => "1001101000000100", 8745 => "1100000011110011", 8746 => "1101111000101100", 8747 => "1111001111111001", 8748 => "0111001111011010", 8749 => "1101101111001001", 8750 => "0011111101111110", 8751 => "0011111110001100", 8752 => "0110010100110010", 8753 => "0010001010010100", 8754 => "0101110001000111", 8755 => "0110010110010000", 8756 => "1100001010101010", 8757 => "1011010110000000", 8758 => "0100111100010111", 8759 => "0011010101100011", 8760 => "1000010110011001", 8761 => "1101111001000110", 8762 => "0111001010000001", 8763 => "1111110011011100", 8764 => "0011000010000000", 8765 => "0010000000011010", 8766 => "1101000101111000", 8767 => "0011110111001000", 8768 => "0001100110100000", 8769 => "0110010001100110", 8770 => "1111110100000000", 8771 => "1000110101011100", 8772 => "0011000101001001", 8773 => "0011111110011010", 8774 => "0100101001100010", 8775 => "0010110001111010", 8776 => "1111001100011010", 8777 => "0010001110000010", 8778 => "1101000000000111", 8779 => "0011101101001111", 8780 => "1011111001001001", 8781 => "1011101010101001", 8782 => "1011001101010101", 8783 => "0010010110100001", 8784 => "1110000110001001", 8785 => "1010110110011011", 8786 => "0010111101100001", 8787 => "1010100111001110", 8788 => "1100010100101100", 8789 => "1011110100110110", 8790 => "1001111101100111", 8791 => "0101100011110000", 8792 => "1110011000100111", 8793 => "0011111111001111", 8794 => "0100001101111011", 8795 => "1011001101000100", 8796 => "0101011101110000", 8797 => "0010001101101000", 8798 => "1101000100010010", 8799 => "0110110001011101", 8800 => "1000101011011100", 8801 => "0100110011111011", 8802 => "0000101001100010", 8803 => "0010101111111110", 8804 => "0010010001011001", 8805 => "1100110011100101", 8806 => "1001000010110001", 8807 => "0000101000101010", 8808 => "0010001001100100", 8809 => "1101010110111100", 8810 => "0111100111110110", 8811 => "0011000010100111", 8812 => "0001111010000101", 8813 => "1110111011100100", 8814 => "1111101010011011", 8815 => "1001110000111000", 8816 => "1010011111101001", 8817 => "0100101000100111", 8818 => "1110100011001111", 8819 => "1000110010011011", 8820 => "0010111000101000", 8821 => "1010101010010111", 8822 => "1000010111001101", 8823 => "0101101001110100", 8824 => "0100000111100101", 8825 => "1110011010101001", 8826 => "0000101100111010", 8827 => "0000001001001101", 8828 => "0100110111001000", 8829 => "1101101011111110", 8830 => "0011010011010111", 8831 => "1000111010111001", 8832 => "1010001001010001", 8833 => "1001100101100000", 8834 => "0001111111011100", 8835 => "1111101011101100", 8836 => "1010010110100000", 8837 => "0000110001111111", 8838 => "0011111001010110", 8839 => "0011011110101101", 8840 => "1010101010110110", 8841 => "0010111010010111", 8842 => "0011011001001110", 8843 => "1110010000100111", 8844 => "0101010001100101", 8845 => "1001011100001000", 8846 => "0011110000000000", 8847 => "0010010000110111", 8848 => "0010111111000100", 8849 => "1001001010100110", 8850 => "0100011010110011", 8851 => "0100111110001111", 8852 => "1111010011010110", 8853 => "0001011000100111", 8854 => "1000010100111010", 8855 => "0001010011111001", 8856 => "1101100101010111", 8857 => "1100100110001110", 8858 => "0011101101111111", 8859 => "0110000110100011", 8860 => "0011100011110000", 8861 => "1101110010000001", 8862 => "1000100010001101", 8863 => "0110101011110101", 8864 => "0000101111100010", 8865 => "0110111000110001", 8866 => "0111101100010010", 8867 => "1110000100011010", 8868 => "0001000111000111", 8869 => "1001000010101000", 8870 => "0011100110001110", 8871 => "1111101111001011", 8872 => "0011101000010111", 8873 => "0001101100010111", 8874 => "0001011000100011", 8875 => "1101110011001100", 8876 => "1110111111100011", 8877 => "0111101001101110", 8878 => "0100101010110000", 8879 => "1101000100110001", 8880 => "1110010010001001", 8881 => "0000011010010010", 8882 => "1101100100101000", 8883 => "0111010100010110", 8884 => "1010001110111111", 8885 => "0001001100000100", 8886 => "0111100110110111", 8887 => "0011011101000101", 8888 => "0011000101111001", 8889 => "1100110001111001", 8890 => "0001100110011010", 8891 => "1000100000000101", 8892 => "0110111001100001", 8893 => "1111100101110100", 8894 => "0000110100100010", 8895 => "0110011101010011", 8896 => "0111101011101111", 8897 => "1000001010001010", 8898 => "0100010000100010", 8899 => "1100001010111100", 8900 => "1101001110011100", 8901 => "0110000010010001", 8902 => "0010010000110100", 8903 => "0011011010000101", 8904 => "0110111010010110", 8905 => "0100011011101010", 8906 => "0100001111100111", 8907 => "0000001010000011", 8908 => "0011101101000111", 8909 => "0110010101001100", 8910 => "1111010100000111", 8911 => "1000100010000100", 8912 => "0111010000011110", 8913 => "0010101000010000", 8914 => "1011010111000111", 8915 => "0011101010000011", 8916 => "0101000111100100", 8917 => "1001011111011010", 8918 => "1000111000001110", 8919 => "0000001011100010", 8920 => "1100111100110011", 8921 => "1110000011010100", 8922 => "1111011101111111", 8923 => "0011011011110101", 8924 => "0110110000100000", 8925 => "1010111101100101", 8926 => "1101000111110110", 8927 => "0110100101110001", 8928 => "0110111010100001", 8929 => "1111010010110111", 8930 => "0100000110010001", 8931 => "1101000111000001", 8932 => "1011001100111111", 8933 => "1011100100001001", 8934 => "0100111110100000", 8935 => "0000011111110010", 8936 => "0000001001111100", 8937 => "0110111101110011", 8938 => "1101011100110100", 8939 => "0110101101111111", 8940 => "1000010100100001", 8941 => "0111100000111000", 8942 => "1010100001110010", 8943 => "1110111101001111", 8944 => "1111000111000110", 8945 => "1000000110111100", 8946 => "0111000010100101", 8947 => "0010100100111111", 8948 => "1001011010011100", 8949 => "1000000001100010", 8950 => "0011001000001101", 8951 => "1100101101110110", 8952 => "0111000010111110", 8953 => "0100010000001110", 8954 => "1110010010111101", 8955 => "0100010011111010", 8956 => "1001111011101110", 8957 => "1101000011011000", 8958 => "1111111110000011", 8959 => "1111011111101000", 8960 => "0111101100010101", 8961 => "0000010101110001", 8962 => "1001011011000111", 8963 => "1010110000000100", 8964 => "0000010011001111", 8965 => "1010100001111110", 8966 => "0001010010110000", 8967 => "0001010010100011", 8968 => "0011111111110011", 8969 => "1001111001000000", 8970 => "1010111001110011", 8971 => "0011100110001101", 8972 => "1110010011010001", 8973 => "1000110111101001", 8974 => "0001100101001011", 8975 => "0110000000110111", 8976 => "0100001110010011", 8977 => "1100001100000001", 8978 => "0110011001000100", 8979 => "0011000000000100", 8980 => "1000101100100000", 8981 => "0100111111010000", 8982 => "0011010110000101", 8983 => "0111101010100010", 8984 => "1001011110100011", 8985 => "1100010100101101", 8986 => "1111010100000100", 8987 => "1100101110010000", 8988 => "0100010110011010", 8989 => "1011001010110111", 8990 => "1100000101100100", 8991 => "0001000110100110", 8992 => "0110010010100010", 8993 => "1110000010011011", 8994 => "1000001111011011", 8995 => "0100111111011100", 8996 => "1100010110101011", 8997 => "0101001110000001", 8998 => "1000011010101011", 8999 => "1100001010011111", 9000 => "1010000101010101", 9001 => "0001111100100001", 9002 => "0100001001101100", 9003 => "1100111110000111", 9004 => "1101111111100111", 9005 => "1111110001000000", 9006 => "0001010100010011", 9007 => "1010010011111101", 9008 => "1010101100010001", 9009 => "1010000101101110", 9010 => "1100111000111001", 9011 => "0001101111000100", 9012 => "1101001111000011", 9013 => "1101101110101010", 9014 => "0111010011101101", 9015 => "1101101101000110", 9016 => "0001100011001100", 9017 => "1011001011001111", 9018 => "1101111011101010", 9019 => "0111011011010001", 9020 => "1011111100100110", 9021 => "1101000011001010", 9022 => "1000111000101101", 9023 => "1010100010101010", 9024 => "1110110111100110", 9025 => "0100011011011011", 9026 => "0110110000001000", 9027 => "1000111000111010", 9028 => "0110011100011001", 9029 => "1100000100001110", 9030 => "0101110000100110", 9031 => "1001000010000110", 9032 => "0101010000010000", 9033 => "0001100100100101", 9034 => "1110111000000101", 9035 => "0111001001111101", 9036 => "0011110111110111", 9037 => "1100101111100110", 9038 => "0011001111010010", 9039 => "1110011100010100", 9040 => "0100100000010001", 9041 => "1000000100010010", 9042 => "0000100010100101", 9043 => "1111111011000011", 9044 => "0011010101110011", 9045 => "1001011110000001", 9046 => "0011110101000011", 9047 => "0101001101101001", 9048 => "1110001101000010", 9049 => "1101010101100010", 9050 => "0100010001101011", 9051 => "1010000110110010", 9052 => "0010111101101000", 9053 => "1010100000100101", 9054 => "1101001000011001", 9055 => "1000000010101010", 9056 => "0101001100001001", 9057 => "0000011001111000", 9058 => "1111000101111000", 9059 => "0000101000011110", 9060 => "0001010001000010", 9061 => "1000101100100000", 9062 => "1110000001111111", 9063 => "1000111000011101", 9064 => "1001110110001011", 9065 => "1011000010001100", 9066 => "0001100110111001", 9067 => "1010100110000110", 9068 => "0010111111001000", 9069 => "1110101101001110", 9070 => "1111111111010011", 9071 => "0111011101110010", 9072 => "1000011011101100", 9073 => "1001111111100000", 9074 => "0001101100111100", 9075 => "0011110011100011", 9076 => "0001001100000001", 9077 => "1100101000101111", 9078 => "1010010011000001", 9079 => "0000111001101000", 9080 => "1010100110001010", 9081 => "0101011100000110", 9082 => "0010000010110110", 9083 => "1010000100100000", 9084 => "1101111011000001", 9085 => "0010101010010001", 9086 => "0101101101101001", 9087 => "0110100101011111", 9088 => "1000111100111000", 9089 => "1110000000011110", 9090 => "1010100011100001", 9091 => "0010010101011011", 9092 => "1001100000111010", 9093 => "1110011101000101", 9094 => "0000100000100110", 9095 => "0111110010111001", 9096 => "1110100101000110", 9097 => "1110011011101110", 9098 => "0001001101100011", 9099 => "0111101100101101", 9100 => "1100110101011011", 9101 => "0110011110001101", 9102 => "0001010110111000", 9103 => "1011011000111010", 9104 => "1100111101000101", 9105 => "1011111111001001", 9106 => "0111110110001110", 9107 => "1000111110011001", 9108 => "1001011111011000", 9109 => "1010010110000010", 9110 => "0001000110111101", 9111 => "0000000011001001", 9112 => "1100000111010000", 9113 => "1000001100000001", 9114 => "1101011100100100", 9115 => "0001011101101001", 9116 => "0010110100101001", 9117 => "0111011111110100", 9118 => "1101101111110000", 9119 => "0001101110110010", 9120 => "0111011110110101", 9121 => "1001111110001011", 9122 => "0001110011001001", 9123 => "1001001010101110", 9124 => "0000100000000100", 9125 => "1100100010010111", 9126 => "1011100011011010", 9127 => "0100010001001110", 9128 => "0011110001000001", 9129 => "1001011001100111", 9130 => "0011001000000001", 9131 => "0011001111000111", 9132 => "1101111011101010", 9133 => "0010111110000011", 9134 => "1100011010110011", 9135 => "0001110001101100", 9136 => "1100111011001000", 9137 => "1101011011000011", 9138 => "1101110000000011", 9139 => "1100101111001111", 9140 => "0110110001001100", 9141 => "1001111101110101", 9142 => "0010101010001110", 9143 => "0111101000000001", 9144 => "1110110100001010", 9145 => "1100001001101010", 9146 => "1110101110101111", 9147 => "1000101111011010", 9148 => "0101010100010001", 9149 => "0111110001001110", 9150 => "1001100100010111", 9151 => "1000111001101001", 9152 => "1000000111000001", 9153 => "0101111011001011", 9154 => "1010110011101000", 9155 => "1000010100001100", 9156 => "1111000110101111", 9157 => "1101010001101001", 9158 => "0011110100110010", 9159 => "1011000110011000", 9160 => "0111110100110001", 9161 => "1101101000000000", 9162 => "1010010011000000", 9163 => "0010000100010100", 9164 => "0010010110011111", 9165 => "1101100001111000", 9166 => "0110111100011101", 9167 => "0111011101101101", 9168 => "0010001111010000", 9169 => "1100011010100100", 9170 => "0010001110001100", 9171 => "0001110011001111", 9172 => "1100101110001110", 9173 => "1111100010110000", 9174 => "0110011111001110", 9175 => "1010110011010000", 9176 => "0011101101011001", 9177 => "0110110101111100", 9178 => "0101100100110001", 9179 => "1101010110101111", 9180 => "1111011001001011", 9181 => "0001001011011010", 9182 => "0011011100111001", 9183 => "1111010000111001", 9184 => "1101001011010110", 9185 => "0100110000001010", 9186 => "0101100001010101", 9187 => "1010001010011010", 9188 => "0000010111011011", 9189 => "1000010000011100", 9190 => "0010101000000010", 9191 => "1110001101100100", 9192 => "0101111111101011", 9193 => "1101110100010001", 9194 => "1111011100000000", 9195 => "0111101110100100", 9196 => "1001000011111101", 9197 => "1101010111010011", 9198 => "1011001000000001", 9199 => "0111111011000111", 9200 => "0000000101110001", 9201 => "0100010111001111", 9202 => "0010101010011000", 9203 => "0100010110000111", 9204 => "0010011000110100", 9205 => "0001000111000110", 9206 => "0110010001010011", 9207 => "0110011101001010", 9208 => "0101110111001011", 9209 => "1111111000111010", 9210 => "1110111101001101", 9211 => "0111110010010001", 9212 => "1101100111111110", 9213 => "1100001000001000", 9214 => "0101010110000000", 9215 => "0100011001101100", 9216 => "1111001101010111", 9217 => "0100111001000101", 9218 => "1001001110000111", 9219 => "0100100111000101", 9220 => "0100100001100101", 9221 => "1011110111111101", 9222 => "1001100100000001", 9223 => "0101110000000000", 9224 => "0011001011101000", 9225 => "0101001111101111", 9226 => "0100010000011011", 9227 => "1001010100101101", 9228 => "0000101101001100", 9229 => "1101011100001001", 9230 => "1110010000011000", 9231 => "1110001001101100", 9232 => "1110010001110101", 9233 => "1111100010110011", 9234 => "1011011001100001", 9235 => "1011111001001011", 9236 => "0100001110000010", 9237 => "1111010011001100", 9238 => "1110001010111010", 9239 => "1000011110100100", 9240 => "1000110111110101", 9241 => "0100101110100100", 9242 => "1110101110010100", 9243 => "0111101101011001", 9244 => "0011000111101100", 9245 => "1110111100110101", 9246 => "0001101000011111", 9247 => "0011000001101011", 9248 => "0010001001111110", 9249 => "1011011010010111", 9250 => "0001110111011011", 9251 => "1010101101100000", 9252 => "0111110011111111", 9253 => "0001011111110101", 9254 => "1011101100101111", 9255 => "0111100110010111", 9256 => "0110111010001100", 9257 => "0010000101001111", 9258 => "0011111101010000", 9259 => "0100011111000110", 9260 => "0011010011011110", 9261 => "0001100011111000", 9262 => "1111001111000010", 9263 => "0100000000110111", 9264 => "1011011011110011", 9265 => "0101110000111111", 9266 => "0010100101011010", 9267 => "1010100000111111", 9268 => "0100000010111001", 9269 => "0011001100000010", 9270 => "0010010110011111", 9271 => "0010100100010000", 9272 => "1001110100110010", 9273 => "1111000111110100", 9274 => "1111111110010101", 9275 => "0001001100110101", 9276 => "0101010101100010", 9277 => "0010000010110001", 9278 => "0100110000001110", 9279 => "0011001001101011", 9280 => "1110111001011000", 9281 => "1011100000101001", 9282 => "1001010001010001", 9283 => "0011010110111010", 9284 => "0000110001011000", 9285 => "1110011111111100", 9286 => "0010011100100111", 9287 => "0101111010111101", 9288 => "1110100101010011", 9289 => "1010000001011101", 9290 => "0100110100111000", 9291 => "1100110100101010", 9292 => "0010011100010110", 9293 => "0000101101110000", 9294 => "0110011100101110", 9295 => "1000001111110001", 9296 => "1010000100101000", 9297 => "1010110101011000", 9298 => "1011011010100111", 9299 => "1100111100010100", 9300 => "0111000001100111", 9301 => "1111001101110000", 9302 => "0101111111010111", 9303 => "0010000100101000", 9304 => "1101111101000110", 9305 => "1010111101100000", 9306 => "1010001101010111", 9307 => "1110110010100000", 9308 => "1011010011111111", 9309 => "0100000001101101", 9310 => "0011101001110111", 9311 => "1010111000101010", 9312 => "1100111101001110", 9313 => "1001101010111100", 9314 => "0000010010110001", 9315 => "0100001101110000", 9316 => "0001100011011000", 9317 => "0010100111011001", 9318 => "0011000101111010", 9319 => "0111001110110110", 9320 => "1001101010011010", 9321 => "1011010100100011", 9322 => "0100001001011000", 9323 => "0100010000011010", 9324 => "0001101011100011", 9325 => "1100000101011001", 9326 => "0011001000100001", 9327 => "0110110110111001", 9328 => "0011001001000101", 9329 => "0100100001101110", 9330 => "1110101010110010", 9331 => "0000000011001111", 9332 => "0000011110010110", 9333 => "1000111100101001", 9334 => "1001010011101100", 9335 => "1110011011101001", 9336 => "1001101011011001", 9337 => "1011110110001011", 9338 => "0011000110101111", 9339 => "1111111110111010", 9340 => "1101001000110010", 9341 => "1101110000011001", 9342 => "0101001110010001", 9343 => "1100111100011110", 9344 => "1001111100101101", 9345 => "0111011001111110", 9346 => "0111010100001111", 9347 => "0000011000111011", 9348 => "1100110111000100", 9349 => "0000011001110101", 9350 => "1010111111101101", 9351 => "1011101001010101", 9352 => "0011001111010111", 9353 => "1001101101011010", 9354 => "1111010111101101", 9355 => "1001101100101000", 9356 => "0010010000010101", 9357 => "0111111111010110", 9358 => "1101100001100101", 9359 => "0000010111000000", 9360 => "0011001100001001", 9361 => "0011111010100110", 9362 => "1010001011110011", 9363 => "1010111000010010", 9364 => "0110001001111010", 9365 => "1000001011110000", 9366 => "1101111000001110", 9367 => "1101110011110100", 9368 => "0110111000010010", 9369 => "0111000000010010", 9370 => "1000101111101110", 9371 => "1011010110000100", 9372 => "1011111010011101", 9373 => "0000100101001000", 9374 => "0100001111010111", 9375 => "0010111101101101", 9376 => "1000010110111001", 9377 => "1001101011001000", 9378 => "0011111110100010", 9379 => "1100110011010000", 9380 => "0110101101011100", 9381 => "0101110000001000", 9382 => "1000111010111111", 9383 => "0000111101001110", 9384 => "1010111110111011", 9385 => "1110110101101101", 9386 => "1011100110110000", 9387 => "1100101111100100", 9388 => "0011111101010111", 9389 => "1011010001101011", 9390 => "1100010011111000", 9391 => "1010111011011110", 9392 => "1111101000101101", 9393 => "0001100010110111", 9394 => "0111000110101000", 9395 => "0000101111101111", 9396 => "1110011011100011", 9397 => "1001110101101101", 9398 => "0110111010000011", 9399 => "1000010000001111", 9400 => "0110010111110111", 9401 => "1000001011011010", 9402 => "0000110010100000", 9403 => "1011010110011010", 9404 => "0011010001000100", 9405 => "1111110111000010", 9406 => "0101100011001011", 9407 => "1011100101010000", 9408 => "1101101100110000", 9409 => "0001000101100100", 9410 => "0000100110001010", 9411 => "1111010111000101", 9412 => "0000110001011011", 9413 => "0110111000100111", 9414 => "1001011011010110", 9415 => "1001000010010101", 9416 => "1010001000100001", 9417 => "0111001001010110", 9418 => "1100110100011100", 9419 => "1001010100101111", 9420 => "1100101110011111", 9421 => "0110100000000001", 9422 => "0010001100101000", 9423 => "0101100101110111", 9424 => "0001101111011000", 9425 => "1000000001111001", 9426 => "1001011011100100", 9427 => "0011001111000110", 9428 => "1100000110101110", 9429 => "1111001111110010", 9430 => "1111111010000111", 9431 => "0001111101010110", 9432 => "0000010001000111", 9433 => "0001110101101001", 9434 => "0000111001010101", 9435 => "1001010010011000", 9436 => "1011001010101000", 9437 => "0000000000111100", 9438 => "0100000010110011", 9439 => "1010100110101111", 9440 => "1100001100110100", 9441 => "0001111000001111", 9442 => "0111001010001001", 9443 => "0110110100100010", 9444 => "0011000100111001", 9445 => "0010001000100011", 9446 => "1000011100111011", 9447 => "0000000011100000", 9448 => "1011110101100001", 9449 => "1100110100011110", 9450 => "1000010010110010", 9451 => "0000000101011001", 9452 => "1100101011000010", 9453 => "0111101101000101", 9454 => "0000000110001111", 9455 => "0000100101011101", 9456 => "1110010001011001", 9457 => "1100010100111011", 9458 => "0111100010110000", 9459 => "1110000011000011", 9460 => "0110101100111000", 9461 => "0000011000111000", 9462 => "1101001001101110", 9463 => "0100011101100111", 9464 => "0010001100100001", 9465 => "0011110100000100", 9466 => "0110011011000111", 9467 => "1011010010111100", 9468 => "1101101011001011", 9469 => "0010011011000010", 9470 => "0111000101000011", 9471 => "1111111101101110", 9472 => "0100110010100111", 9473 => "1000111000101001", 9474 => "1000000100111101", 9475 => "1111000110010001", 9476 => "1110001110000111", 9477 => "1001100101000000", 9478 => "1100100000011000", 9479 => "1101111100010101", 9480 => "0001001100111110", 9481 => "0000010110000010", 9482 => "1111001001100000", 9483 => "0010001001111101", 9484 => "1010100011101111", 9485 => "1010101000000001", 9486 => "0100101000001111", 9487 => "1111001010011011", 9488 => "0011110100010001", 9489 => "0000100010001110", 9490 => "1011111110010010", 9491 => "0111111000101001", 9492 => "0110101010011000", 9493 => "1011100100011010", 9494 => "1000011101011110", 9495 => "0000111110101000", 9496 => "1101111000011111", 9497 => "1110111110101110", 9498 => "1000110010001111", 9499 => "0111111101100101", 9500 => "0100101010110100", 9501 => "0110011110100001", 9502 => "1101000111110101", 9503 => "1010111111111100", 9504 => "0010010000111100", 9505 => "1000101010101011", 9506 => "1000011001010000", 9507 => "0100110011110000", 9508 => "0110101010001011", 9509 => "1110000001000111", 9510 => "1001011000110110", 9511 => "1010000111111000", 9512 => "0010101101110000", 9513 => "0010001110010101", 9514 => "0011111101110011", 9515 => "1000111000101101", 9516 => "0111011001111111", 9517 => "1100100001010010", 9518 => "0110111011010011", 9519 => "0101000011000101", 9520 => "0111011010100110", 9521 => "0011100000111001", 9522 => "1101010000110000", 9523 => "1101101010011011", 9524 => "1111001111100110", 9525 => "1100111110101011", 9526 => "0000010010101010", 9527 => "1000001000001000", 9528 => "0011001001111010", 9529 => "1111011000111000", 9530 => "1111101111101110", 9531 => "0110100100001111", 9532 => "1010011000110101", 9533 => "0101011100010001", 9534 => "0001110000011101", 9535 => "0001010010101100", 9536 => "1110000011100001", 9537 => "1100000000000000", 9538 => "1001000100101001", 9539 => "0011011110110100", 9540 => "1001010001010111", 9541 => "0000000100100110", 9542 => "1011110101000110", 9543 => "0010000011010011", 9544 => "1001001100110000", 9545 => "1011111000110011", 9546 => "0010011110110000", 9547 => "1011111000001011", 9548 => "1001101010100110", 9549 => "1011111011001010", 9550 => "0010010100010100", 9551 => "0001110100001011", 9552 => "0101000000011111", 9553 => "1011111100000010", 9554 => "0001101001011001", 9555 => "1101000000010001", 9556 => "0011010001110010", 9557 => "1010110110000010", 9558 => "0001100001011000", 9559 => "1110010011010101", 9560 => "1101011101100101", 9561 => "1010001111011011", 9562 => "1000000111111001", 9563 => "0011001000011011", 9564 => "0110110001011001", 9565 => "0110000100010011", 9566 => "1010010110101110", 9567 => "1011111100111001", 9568 => "1100011010110011", 9569 => "1010111010100011", 9570 => "1110101010000001", 9571 => "0100011110000000", 9572 => "0001001100001111", 9573 => "1010111000011110", 9574 => "1110100111111111", 9575 => "1101000101000101", 9576 => "0100001000000111", 9577 => "0110000101000111", 9578 => "0001000010010100", 9579 => "1100111111100101", 9580 => "1110001010111100", 9581 => "1101111111001010", 9582 => "0001111001101001", 9583 => "1101111100000100", 9584 => "0110001011100010", 9585 => "0010001100111101", 9586 => "1010000111101001", 9587 => "1101101110111010", 9588 => "1001101010100011", 9589 => "1001100000111111", 9590 => "1110001101011010", 9591 => "0010111110100011", 9592 => "1111010011011110", 9593 => "0011111010001001", 9594 => "0101000001010101", 9595 => "0000010100011010", 9596 => "1010000101111001", 9597 => "1001101011100000", 9598 => "0011101001000001", 9599 => "1110111011010011", 9600 => "1100011010001000", 9601 => "1011100101010000", 9602 => "1100010000101011", 9603 => "0010000011101110", 9604 => "1110101101101000", 9605 => "0000010011001110", 9606 => "1001000111100010", 9607 => "1000101110101100", 9608 => "0101101001010010", 9609 => "1010000111010100", 9610 => "0110100000001100", 9611 => "1101000001010111", 9612 => "1110011100010110", 9613 => "0100111010011110", 9614 => "0010000111001000", 9615 => "1111111111000000", 9616 => "1001100000010001", 9617 => "1010100011100001", 9618 => "0000101100010111", 9619 => "0101110000001001", 9620 => "0011010011111101", 9621 => "1111011110100100", 9622 => "1100110111000000", 9623 => "1100010000010010", 9624 => "1111110010101110", 9625 => "1110101100001111", 9626 => "0111111100101001", 9627 => "1111001011111000", 9628 => "0111011010010011", 9629 => "1010111010100110", 9630 => "0100111011010001", 9631 => "1010001101000100", 9632 => "1010100110110011", 9633 => "0100111101001111", 9634 => "1111011111111010", 9635 => "0000001000011111", 9636 => "1100101110101110", 9637 => "0110110110000100", 9638 => "0011111101101001", 9639 => "1000110010101001", 9640 => "1110001011000100", 9641 => "0101111001100011", 9642 => "1111111111010110", 9643 => "1001101011110110", 9644 => "1100001110110101", 9645 => "0010111000110101", 9646 => "0110100110000100", 9647 => "1101100111100100", 9648 => "1000000010111010", 9649 => "0101000100010111", 9650 => "0000101011111100", 9651 => "1110000110000110", 9652 => "1011000000001000", 9653 => "0110001000001110", 9654 => "1100110110001111", 9655 => "0111000101011010", 9656 => "1000110011001010", 9657 => "0100110010001000", 9658 => "1011011110101111", 9659 => "0111010111001100", 9660 => "0100110011001010", 9661 => "0010100001000111", 9662 => "0100001110001110", 9663 => "1111011000100010", 9664 => "1110011111010110", 9665 => "1011110111100011", 9666 => "1001111000100101", 9667 => "1000011100111001", 9668 => "0100001011010010", 9669 => "0010011000000001", 9670 => "0101010101010100", 9671 => "0011110001101001", 9672 => "1000101111000110", 9673 => "0001100000010011", 9674 => "0000110011100101", 9675 => "0000011001111110", 9676 => "1111011110001000", 9677 => "0111110000100001", 9678 => "0110001110010010", 9679 => "1001101101110011", 9680 => "0000001011111101", 9681 => "1111101011001010", 9682 => "0101010011000101", 9683 => "0011100101011001", 9684 => "1010010000011100", 9685 => "0010111110010111", 9686 => "0110110011111101", 9687 => "1001011101010010", 9688 => "0001010011110101", 9689 => "0110000101011101", 9690 => "0000001101010110", 9691 => "1001101110110010", 9692 => "1000001001111100", 9693 => "1101001000011101", 9694 => "0101011101110011", 9695 => "1111101011100101", 9696 => "1111001101000010", 9697 => "1011111101100001", 9698 => "1010001101011100", 9699 => "1001111000000101", 9700 => "1010010001000110", 9701 => "0110110111011110", 9702 => "1011101000010110", 9703 => "0110100010010000", 9704 => "1000010011101111", 9705 => "0011010110101100", 9706 => "0001100110110110", 9707 => "0001000110001010", 9708 => "0110010100101011", 9709 => "0101000111011101", 9710 => "1100001101011000", 9711 => "1111101111110110", 9712 => "0111100001000101", 9713 => "0000111111110001", 9714 => "0101110010011110", 9715 => "1111001001100111", 9716 => "1010100010000010", 9717 => "1111110010010101", 9718 => "0101110001011001", 9719 => "1101001001101010", 9720 => "0111110011010100", 9721 => "1001011000000001", 9722 => "0111100110001100", 9723 => "1010010100110011", 9724 => "0010111101101001", 9725 => "1110000011100001", 9726 => "1110011001110110", 9727 => "0000010100101111", 9728 => "1010101000110100", 9729 => "0101010111000100", 9730 => "1111010001001101", 9731 => "1101010011111010", 9732 => "1101101100110011", 9733 => "0011101101001000", 9734 => "0011010000011111", 9735 => "0100001111001111", 9736 => "0101001110100011", 9737 => "0010000000011010", 9738 => "0100001000001101", 9739 => "1011010000010001", 9740 => "1110010111001100", 9741 => "1100010001111010", 9742 => "1000001101101110", 9743 => "1101011111010100", 9744 => "1011100001110100", 9745 => "1010000100100001", 9746 => "0001001001111010", 9747 => "0011011001001010", 9748 => "0110101001101111", 9749 => "0011011110101011", 9750 => "1000100100111110", 9751 => "1010110010010011", 9752 => "1010000000101101", 9753 => "0101110000111111", 9754 => "0101001000101110", 9755 => "1001110111100011", 9756 => "0101011001011110", 9757 => "0101110110100011", 9758 => "0000111110110010", 9759 => "1011000111100111", 9760 => "1010010110001101", 9761 => "1001001110110010", 9762 => "0100111101001100", 9763 => "0010100100000111", 9764 => "1000100101000000", 9765 => "1001001100100101", 9766 => "0100111110011000", 9767 => "0001110001001110", 9768 => "1011100111011010", 9769 => "1010100100000010", 9770 => "0111111100111000", 9771 => "1010001010100100", 9772 => "0001000111010100", 9773 => "0100110001011110", 9774 => "1111010111111001", 9775 => "1011000001001110", 9776 => "0110011101010010", 9777 => "1001101011010000", 9778 => "1100010100101011", 9779 => "1110000110000111", 9780 => "0110011100011111", 9781 => "1010010110110101", 9782 => "0011001111001100", 9783 => "1100110110000001", 9784 => "0001110110000010", 9785 => "0111011000010100", 9786 => "0101110110011101", 9787 => "0101011101010000", 9788 => "1000101010110000", 9789 => "1101001010010110", 9790 => "1111101011111100", 9791 => "0101010100011100", 9792 => "0111101110011101", 9793 => "0001010011110011", 9794 => "0010001101111101", 9795 => "1001111111110110", 9796 => "1111011001100101", 9797 => "1010101110111110", 9798 => "1001111001110110", 9799 => "1101111111010101", 9800 => "1001110001101111", 9801 => "1001111001110100", 9802 => "1110100110001000", 9803 => "0101000111110111", 9804 => "0011000000111111", 9805 => "1111010101101011", 9806 => "1110111000101010", 9807 => "0010100010010011", 9808 => "0111000000001000", 9809 => "0010100111000111", 9810 => "0110000000010000", 9811 => "0111100100110001", 9812 => "1010011101010101", 9813 => "1111010000100010", 9814 => "1001001001111101", 9815 => "0011101100001100", 9816 => "1100101010011110", 9817 => "1011010110111101", 9818 => "0101110000011100", 9819 => "1111110001111010", 9820 => "0100110010110110", 9821 => "1010010011011111", 9822 => "1101110000001001", 9823 => "1011110010100101", 9824 => "1100010100101010", 9825 => "0101011111110000", 9826 => "1101011101110000", 9827 => "1010111101110111", 9828 => "0111001000000000", 9829 => "0100011100111100", 9830 => "1111101001001011", 9831 => "1110101111010110", 9832 => "0001110110011001", 9833 => "0010000101000100", 9834 => "0000001111100111", 9835 => "1110110000110000", 9836 => "0011000000001000", 9837 => "1011110110101001", 9838 => "0110010111011101", 9839 => "1011000111001011", 9840 => "1011101011010001", 9841 => "1100111010110000", 9842 => "1010000110011011", 9843 => "0010100001000001", 9844 => "0101110001011011", 9845 => "1010000100100101", 9846 => "1110000011101001", 9847 => "0101100111000010", 9848 => "0000001000001001", 9849 => "0011111110110010", 9850 => "0101000101000100", 9851 => "0000101100001101", 9852 => "1001011101110101", 9853 => "1001001000000000", 9854 => "1001001011101001", 9855 => "1001101101000100", 9856 => "0101100110000010", 9857 => "1000001000011101", 9858 => "0001001000001010", 9859 => "1100110111110100", 9860 => "0111011000010001", 9861 => "0011101111000100", 9862 => "1001011100110101", 9863 => "0111011111110111", 9864 => "0011001100111111", 9865 => "0111010001010011", 9866 => "0000010110011011", 9867 => "1100110111010110", 9868 => "1001011010001110", 9869 => "1011110011010000", 9870 => "0111110001100111", 9871 => "1010101011010001", 9872 => "1101110011000110", 9873 => "0101010010001111", 9874 => "0111111011110000", 9875 => "0100101101101111", 9876 => "1000101110001101", 9877 => "1000100011110110", 9878 => "0101000000011111", 9879 => "1011000011110100", 9880 => "0111101010010010", 9881 => "1000110100101010", 9882 => "1110101110110101", 9883 => "0000100101000010", 9884 => "1000101111010100", 9885 => "0110101001111100", 9886 => "1110101111010011", 9887 => "1001011000000001", 9888 => "0100011000101010", 9889 => "0101001011110000", 9890 => "0001010001011010", 9891 => "1001101111101111", 9892 => "1110011000101000", 9893 => "0010000101001001", 9894 => "0101001100110010", 9895 => "0001111011110101", 9896 => "0110001001101001", 9897 => "1000001111111101", 9898 => "1111000111010110", 9899 => "0110101110011110", 9900 => "0101100010110101", 9901 => "0101011100001001", 9902 => "0011111010011001", 9903 => "0110011101010000", 9904 => "1010001001101101", 9905 => "1101001001010001", 9906 => "1010010001010111", 9907 => "0011111101010010", 9908 => "0100011111000110", 9909 => "1001110101111000", 9910 => "0101001100101011", 9911 => "1100111101000111", 9912 => "0110111100101111", 9913 => "1110001111011000", 9914 => "1001110011011110", 9915 => "0001000011010010", 9916 => "0010010101110001", 9917 => "1000001001101111", 9918 => "1111100000111000", 9919 => "0100011110011000", 9920 => "1001111110101100", 9921 => "0110110100000101", 9922 => "0101010000000110", 9923 => "0111110000010011", 9924 => "1001111001010111", 9925 => "1110101101111010", 9926 => "0000011000110001", 9927 => "0010001000101101", 9928 => "1111111011010100", 9929 => "1001110101110011", 9930 => "1111001111101010", 9931 => "1101011111000101", 9932 => "0011101101101011", 9933 => "0111110110000100", 9934 => "0101010101000001", 9935 => "1111010110001100", 9936 => "0011010000010111", 9937 => "1000100000001110", 9938 => "1100011000000111", 9939 => "0110000111100110", 9940 => "1010100001001100", 9941 => "1101010001000011", 9942 => "1100110100001011", 9943 => "1101101000000110", 9944 => "1100101000001101", 9945 => "0011010010100100", 9946 => "0111011111111001", 9947 => "0010010000101100", 9948 => "1100110010111010", 9949 => "0010111000100010", 9950 => "1110111000010000", 9951 => "1110111001111111", 9952 => "0110110110010010", 9953 => "1100011111011000", 9954 => "0111100100101101", 9955 => "0000110100000000", 9956 => "0100100110000111", 9957 => "0011010111000010", 9958 => "0101010001110011", 9959 => "1010110111100000", 9960 => "0111100000010100", 9961 => "0110100010111100", 9962 => "0010101001010111", 9963 => "1101010110010100", 9964 => "1011110000000110", 9965 => "1011100100010110", 9966 => "0100001011000101", 9967 => "1011100000010001", 9968 => "1111000011001111", 9969 => "1100000111011000", 9970 => "1010110100000000", 9971 => "0011010000100111", 9972 => "0011101011110110", 9973 => "0000001000111010", 9974 => "1010101011100110", 9975 => "0011110010000111", 9976 => "0110101101011010", 9977 => "1011001001101101", 9978 => "1001000010001000", 9979 => "0010001001111011", 9980 => "0110110111000000", 9981 => "1101111011111111", 9982 => "1110100110100110", 9983 => "0110010111011101", 9984 => "0001111110100101", 9985 => "1110110011111101", 9986 => "1011000011010101", 9987 => "1101101001110100", 9988 => "1101011111111010", 9989 => "1111101101111100", 9990 => "1000110010001110", 9991 => "1010001001001100", 9992 => "1001111001011111", 9993 => "1001100110000100", 9994 => "1101001010110101", 9995 => "0100100000001011", 9996 => "0010101000011000", 9997 => "1011000100011111", 9998 => "1100101000001000", 9999 => "0011101000001010", 10000 => "1011100101110110", 10001 => "1100111110110010", 10002 => "1101100110000011", 10003 => "0011000101000001", 10004 => "1100011100011110", 10005 => "0001010111011011", 10006 => "1010001011011001", 10007 => "0100001001001101", 10008 => "0001111100110100", 10009 => "1000101110111011", 10010 => "0110010100011000", 10011 => "0000000100001001", 10012 => "1100111001001001", 10013 => "1000101101000110", 10014 => "1110000100111110", 10015 => "1000011101011001", 10016 => "0011100111010100", 10017 => "1101111110011000", 10018 => "0010011100011111", 10019 => "1011110100110110", 10020 => "0101100100011111", 10021 => "1101111000101010", 10022 => "0100010000110100", 10023 => "0100100100110101", 10024 => "1100011001000010", 10025 => "0101011101100101", 10026 => "0101100000101110", 10027 => "0101101011110010", 10028 => "1011101011101001", 10029 => "1010000000011000", 10030 => "1010111111100101", 10031 => "0111001101100010", 10032 => "0001011000001000", 10033 => "0000111100000100", 10034 => "0001110010101000", 10035 => "1110101101110000", 10036 => "1001111110100010", 10037 => "1110100110010110", 10038 => "1000011000010011", 10039 => "0101100111000011", 10040 => "0110011001100001", 10041 => "1110101100111111", 10042 => "0010110000001010", 10043 => "1110110101101110", 10044 => "1100100001001001", 10045 => "0011101111011101", 10046 => "0011001101101010", 10047 => "1101110011011100", 10048 => "0111110010011000", 10049 => "1100001110110000", 10050 => "0010010011000001", 10051 => "1011111111100101", 10052 => "0010101100101010", 10053 => "1011101000110101", 10054 => "0100011111111011", 10055 => "0100101111101011", 10056 => "0010001000011000", 10057 => "1010001110110100", 10058 => "0111100100010010", 10059 => "1100000100010111", 10060 => "1101101110110110", 10061 => "0010100010001111", 10062 => "1101001101001100", 10063 => "1000001101110110", 10064 => "0100011101010000", 10065 => "0011101110110111", 10066 => "0001110100011011", 10067 => "0111100110001011", 10068 => "0110000010100101", 10069 => "1000000100000001", 10070 => "0011000000101110", 10071 => "0011101110111110", 10072 => "1101110110100100", 10073 => "0101001010110101", 10074 => "1000110101010110", 10075 => "1111000110000101", 10076 => "1000001011110011", 10077 => "1101011001101101", 10078 => "1010011100111110", 10079 => "0000000110111111", 10080 => "0001100010111010", 10081 => "0010100010101011", 10082 => "0011011011111011", 10083 => "0110111100001000", 10084 => "0000001011011010", 10085 => "0011000000100000", 10086 => "1111010100110010", 10087 => "1011011011011010", 10088 => "0011111000011010", 10089 => "1000001101101100", 10090 => "0110011101001111", 10091 => "1011010101110000", 10092 => "0000011100011001", 10093 => "1011101001001001", 10094 => "0000110111110010", 10095 => "1111101001001101", 10096 => "0111001111101000", 10097 => "0101100100011000", 10098 => "0010011100111000", 10099 => "0011001001000001", 10100 => "1000000011001001", 10101 => "0100001001001100", 10102 => "0100001010110100", 10103 => "1110111110110100", 10104 => "0101010010111111", 10105 => "1010101001110001", 10106 => "0101111111101101", 10107 => "0010110101110111", 10108 => "1101111000010000", 10109 => "0101101011100111", 10110 => "0110010000010010", 10111 => "0101100101001001", 10112 => "0100000000010000", 10113 => "1001100111010001", 10114 => "1011011011100110", 10115 => "0010011110001100", 10116 => "1101111001010101", 10117 => "1000010101111011", 10118 => "1001010101111101", 10119 => "0000000011000110", 10120 => "0011101011010111", 10121 => "1011101011101010", 10122 => "1000100110000100", 10123 => "0001100111100111", 10124 => "1100110100101101", 10125 => "1000111100101011", 10126 => "0101010001001100", 10127 => "0101101011011000", 10128 => "0110110101001100", 10129 => "1011010110111110", 10130 => "1010010001110011", 10131 => "1100011111111001", 10132 => "0100010010010010", 10133 => "1100011110111110", 10134 => "1001000000111110", 10135 => "0111011101001011", 10136 => "0010001101001000", 10137 => "0010110101000000", 10138 => "1110101001000001", 10139 => "1000101001000111", 10140 => "0110101000011101", 10141 => "0010010001101011", 10142 => "1100110000101011", 10143 => "0000001101110011", 10144 => "1011010111000011", 10145 => "1111111000101101", 10146 => "0101110011010010", 10147 => "0100111110111001", 10148 => "1101111001111001", 10149 => "1001111001000010", 10150 => "0100100000010111", 10151 => "0111000000011010", 10152 => "1001000110011001", 10153 => "1000100110010101", 10154 => "1101011011110100", 10155 => "0100110010111111", 10156 => "0000111000100010", 10157 => "0000001100101101", 10158 => "0111010110111010", 10159 => "0101001010101101", 10160 => "0101101101100011", 10161 => "1011110101110111", 10162 => "0011010001111010", 10163 => "1011000111110110", 10164 => "1010101110010100", 10165 => "0011000111000111", 10166 => "0110101101111110", 10167 => "0110101010010001", 10168 => "0100100101110011", 10169 => "0001000100110101", 10170 => "1100001000100110", 10171 => "0000110101111000", 10172 => "1001101011011111", 10173 => "0101110000000101", 10174 => "1111001001111011", 10175 => "0001010001000110", 10176 => "1010111110100010", 10177 => "0110011111100100", 10178 => "0011101001000111", 10179 => "0101011100101100", 10180 => "0010100011011011", 10181 => "1100110100100110", 10182 => "0100110101010110", 10183 => "0010100100000011", 10184 => "1110011100011011", 10185 => "1000001101001001", 10186 => "0101110101000101", 10187 => "1001011110000100", 10188 => "0000111100111010", 10189 => "1001000101010011", 10190 => "0010101100110111", 10191 => "1001111000000110", 10192 => "0001010100010011", 10193 => "1101101011111000", 10194 => "0011100011010010", 10195 => "0111111010001010", 10196 => "0011111110010100", 10197 => "0010000011000101", 10198 => "1101100100001000", 10199 => "1001001001010110", 10200 => "0111110111010111", 10201 => "1010111100010000", 10202 => "1010111000110010", 10203 => "0000010010000000", 10204 => "0000110000001111", 10205 => "0111110011111100", 10206 => "1010000111011110", 10207 => "1100001101100000", 10208 => "0011010111001100", 10209 => "0010000110001011", 10210 => "0000001001101100", 10211 => "1010011110000100", 10212 => "1010100010110110", 10213 => "1010101000101010", 10214 => "1000101100010101", 10215 => "1111010000110000", 10216 => "0110111001011000", 10217 => "1010110000111100", 10218 => "1001101010111110", 10219 => "1100101110110000", 10220 => "1011001100100010", 10221 => "1001000101000010", 10222 => "0100010101001001", 10223 => "0111101011110000", 10224 => "0101000100010101", 10225 => "1111001000101110", 10226 => "1000010010111101", 10227 => "0111010000010011", 10228 => "0101001001100000", 10229 => "1000010101011110", 10230 => "1101011001011011", 10231 => "0100001100101001", 10232 => "1000001100110100", 10233 => "0001010110111001", 10234 => "0110010010100111", 10235 => "0110001001001111", 10236 => "1011011111110110", 10237 => "1111001110110110", 10238 => "0010000011000001", 10239 => "1010001000000100", 10240 => "0111000011111111", 10241 => "1010100000110010", 10242 => "0000001001111001", 10243 => "0101101100011111", 10244 => "1101010011011011", 10245 => "0011110000100010", 10246 => "0100010111000100", 10247 => "0110000100010100", 10248 => "0111111110011011", 10249 => "1001001011001010", 10250 => "1101000101101101", 10251 => "1100001011011011", 10252 => "1101111111100111", 10253 => "0010000100010001", 10254 => "1111101011100110", 10255 => "1101100111011011", 10256 => "1111100100000101", 10257 => "0100001000111110", 10258 => "1101110111001011", 10259 => "1011001001000010", 10260 => "1100100101000111", 10261 => "0001110110010110", 10262 => "1001001000011101", 10263 => "1010101011010011", 10264 => "0000110100111111", 10265 => "0001100000010110", 10266 => "1110100110011000", 10267 => "1110101101011011", 10268 => "1110101000110101", 10269 => "0011100001110011", 10270 => "0100001110000011", 10271 => "0110001110000100", 10272 => "1001011000010000", 10273 => "1011101011111111", 10274 => "1111001111101100", 10275 => "1001011101110001", 10276 => "0000010001111001", 10277 => "1010011001101010", 10278 => "1101100101111011", 10279 => "1100110101001111", 10280 => "0011100011001100", 10281 => "0100111000100100", 10282 => "0111000111011011", 10283 => "1000000100111101", 10284 => "1111010010010111", 10285 => "1111100101111001", 10286 => "0110011101111001", 10287 => "0010101100011000", 10288 => "1111010010110111", 10289 => "0001100111000011", 10290 => "0001001101100101", 10291 => "0010000000010000", 10292 => "1001111111001001", 10293 => "0011111001010011", 10294 => "1100101101111111", 10295 => "1110010000010010", 10296 => "0010010101010111", 10297 => "0010111001100100", 10298 => "0001110110000100", 10299 => "1001111000100001", 10300 => "1100010000001010", 10301 => "0111100110011100", 10302 => "0111010011110100", 10303 => "0111010100110101", 10304 => "1110001100010110", 10305 => "1100000010000111", 10306 => "0101110100010101", 10307 => "1011001100011101", 10308 => "1100001110010011", 10309 => "1110100111100100", 10310 => "0011101101000100", 10311 => "1111111111111000", 10312 => "0100000111111011", 10313 => "1110001011101110", 10314 => "1010110101011001", 10315 => "0011111010011101", 10316 => "1000010100000001", 10317 => "0101010001110111", 10318 => "0110011010010010", 10319 => "0011101110010101", 10320 => "1101110111111000", 10321 => "0011110100101001", 10322 => "1010001100000011", 10323 => "0010100010101100", 10324 => "0011110111001011", 10325 => "1001010011010001", 10326 => "1010100011001101", 10327 => "1110110000010000", 10328 => "0001101010111101", 10329 => "1010010000001011", 10330 => "0111001011111010", 10331 => "0010011001101101", 10332 => "0111110100110101", 10333 => "1000100011001010", 10334 => "1001111001111101", 10335 => "0111101110111101", 10336 => "1100000000100101", 10337 => "1001001011001100", 10338 => "1010100101010101", 10339 => "1100100010100100", 10340 => "1100110000110001", 10341 => "0000100101011001", 10342 => "0111110101110010", 10343 => "1100101100001010", 10344 => "1010111010010100", 10345 => "1010111010111110", 10346 => "0100111100111101", 10347 => "0000101010010100", 10348 => "0111011100100110", 10349 => "1010100111011011", 10350 => "1011101100001001", 10351 => "0000011001010010", 10352 => "0110111010110110", 10353 => "1001100111101110", 10354 => "0000110000110000", 10355 => "1011100100001010", 10356 => "0001101001010110", 10357 => "1001110110110101", 10358 => "0111110010000111", 10359 => "1111101100011011", 10360 => "1011011111100101", 10361 => "0001001111100000", 10362 => "0110100010110110", 10363 => "1100110110001011", 10364 => "0110001000111111", 10365 => "0011000001101100", 10366 => "1001001100111111", 10367 => "0001000110001010", 10368 => "1010101101011101", 10369 => "0110100110110100", 10370 => "1011011001001101", 10371 => "0011110111000111", 10372 => "0001000110010100", 10373 => "0000111110110110", 10374 => "0101101010100100", 10375 => "1001000100100111", 10376 => "1000000001100111", 10377 => "0101011110001101", 10378 => "0000101001011100", 10379 => "0110001010101011", 10380 => "1110011010011111", 10381 => "1101010100100101", 10382 => "0110100111010010", 10383 => "0101011010011110", 10384 => "0110101100110101", 10385 => "1101110101000100", 10386 => "0101010101010111", 10387 => "1010101000111001", 10388 => "1100001110001111", 10389 => "0111000101001000", 10390 => "0001110100001001", 10391 => "1001001111111001", 10392 => "1110100010100100", 10393 => "1101100100101100", 10394 => "1011010101100001", 10395 => "0111011000111110", 10396 => "0011001110001101", 10397 => "1110001100000010", 10398 => "0001100110000110", 10399 => "1111110110011110", 10400 => "0110000111010011", 10401 => "1001010000100001", 10402 => "1100110111011111", 10403 => "1000001011001010", 10404 => "1110111010011101", 10405 => "1001000110010101", 10406 => "1100110100011010", 10407 => "1110110100011010", 10408 => "1010100111001000", 10409 => "1011101010000001", 10410 => "0100111110101010", 10411 => "1111000101101100", 10412 => "1011001000001001", 10413 => "0110111001010000", 10414 => "1011001101001100", 10415 => "1101000000100101", 10416 => "1100111100001101", 10417 => "1111010111001001", 10418 => "1110001100000000", 10419 => "0100101110110100", 10420 => "1100001101011110", 10421 => "0100100100000111", 10422 => "0001001010000000", 10423 => "0100010110110000", 10424 => "0010110010011101", 10425 => "1101110011001110", 10426 => "0101011110111010", 10427 => "0010111111100111", 10428 => "0101010001111111", 10429 => "1110011100111010", 10430 => "1110111110101001", 10431 => "0010110100101000", 10432 => "1001011010010110", 10433 => "0111101111101110", 10434 => "0100001010011001", 10435 => "1001110010111110", 10436 => "1001100100011010", 10437 => "0010010011101111", 10438 => "0011100111001011", 10439 => "1001100010101110", 10440 => "0010110000110110", 10441 => "1111100001000110", 10442 => "0110100010110100", 10443 => "0000010000001110", 10444 => "1101110010100011", 10445 => "0001000000010000", 10446 => "1110000110111110", 10447 => "1101100010101011", 10448 => "0100101011010110", 10449 => "0101100011111011", 10450 => "1000011111110000", 10451 => "0001001000110101", 10452 => "1100111001001001", 10453 => "0111010111110011", 10454 => "0010000100011111", 10455 => "0100100010010001", 10456 => "0000001100111011", 10457 => "1101110100000111", 10458 => "0101110001110100", 10459 => "1111000111101001", 10460 => "0000110101111010", 10461 => "0110101111100110", 10462 => "1101100111111100", 10463 => "0001101000010110", 10464 => "1010111011110001", 10465 => "1010111110100010", 10466 => "0000011011001010", 10467 => "0110101001111110", 10468 => "0010001100101010", 10469 => "0111100110000001", 10470 => "1101011110101001", 10471 => "0011111111010000", 10472 => "0010011011000100", 10473 => "1101000010110111", 10474 => "0111111101010110", 10475 => "1000100010111101", 10476 => "1010011010101110", 10477 => "1110000010010011", 10478 => "0011110010100110", 10479 => "0010100100010011", 10480 => "1101000100000110", 10481 => "1110100011110100", 10482 => "0110110010100100", 10483 => "0110010100010000", 10484 => "0110101101010110", 10485 => "0000001111011000", 10486 => "0010000101100010", 10487 => "0101100000000100", 10488 => "0101000110111000", 10489 => "1111101110011111", 10490 => "1011101000101011", 10491 => "0111110010101000", 10492 => "0000001100101010", 10493 => "1100100000101011", 10494 => "1000101000000000", 10495 => "1110111111111101", 10496 => "1101010111110100", 10497 => "0111010000100100", 10498 => "0011111010000010", 10499 => "0000011001010110", 10500 => "1011100010110101", 10501 => "0110110000111110", 10502 => "0101111101010101", 10503 => "0100101001000001", 10504 => "1100000010110000", 10505 => "1011001011001000", 10506 => "0010101100110110", 10507 => "1100100111001110", 10508 => "1011011001010000", 10509 => "0011000010100101", 10510 => "0010100010110011", 10511 => "0110011001011010", 10512 => "1101111010101011", 10513 => "0100011011010100", 10514 => "1110100001110001", 10515 => "1110000100011011", 10516 => "1001011001001101", 10517 => "1010101001010011", 10518 => "1110001011001001", 10519 => "1010100110001100", 10520 => "1100000110001011", 10521 => "0000010011011101", 10522 => "1101010110011111", 10523 => "1011101100000001", 10524 => "0000110000111000", 10525 => "0000101010110101", 10526 => "1101100100101011", 10527 => "1100110000010100", 10528 => "0000010100100100", 10529 => "1000111010001100", 10530 => "1110111101011011", 10531 => "1101111111001011", 10532 => "1101111101010111", 10533 => "1110000010000011", 10534 => "1011011101001110", 10535 => "0101000010011011", 10536 => "1110011001011100", 10537 => "0111100100101110", 10538 => "1110010011000000", 10539 => "0000001010010011", 10540 => "1010011110000111", 10541 => "1011001000100100", 10542 => "1011010101110010", 10543 => "1110101000010011", 10544 => "0101100011010011", 10545 => "1011001101101001", 10546 => "1100111111001001", 10547 => "0111101010101110", 10548 => "1000010010110000", 10549 => "0001101100110100", 10550 => "0011000111100100", 10551 => "1000110101111000", 10552 => "0010011101100110", 10553 => "1000101000001000", 10554 => "0110100100011011", 10555 => "1000010110100110", 10556 => "1001101001111011", 10557 => "0101011000010100", 10558 => "1100000111000000", 10559 => "1010100010101001", 10560 => "0110011101111101", 10561 => "1000111111101010", 10562 => "1011011111011100", 10563 => "1110101001010110", 10564 => "1101101011110111", 10565 => "1000111101110100", 10566 => "0001000101101001", 10567 => "0101111000101011", 10568 => "0000100111011101", 10569 => "0001111010010101", 10570 => "0010011110101001", 10571 => "0001110101100000", 10572 => "0011011000000111", 10573 => "1010100100001011", 10574 => "1101010101000001", 10575 => "0001001010111111", 10576 => "0011100010001001", 10577 => "0001000101111111", 10578 => "1001011010010111", 10579 => "1011100110010011", 10580 => "0000011101011000", 10581 => "0111100110000010", 10582 => "1100111111001101", 10583 => "1000000111101100", 10584 => "0101101011010010", 10585 => "1101100111001110", 10586 => "0100010101111111", 10587 => "1110101110111100", 10588 => "1111110101011110", 10589 => "0011101011111001", 10590 => "1100100110010100", 10591 => "0101101101101011", 10592 => "0010110100110011", 10593 => "0110111111111011", 10594 => "1100101000100000", 10595 => "0000001010000000", 10596 => "1111011100110111", 10597 => "1001001110001001", 10598 => "0010001111000110", 10599 => "0100011000101111", 10600 => "0011111101010000", 10601 => "1010001111011101", 10602 => "0010010111010111", 10603 => "1010000100100001", 10604 => "0111100000001001", 10605 => "0011010011101000", 10606 => "1000111011110100", 10607 => "1111010110000000", 10608 => "1011000100010100", 10609 => "1000101000110111", 10610 => "0011011100001100", 10611 => "1110101101000000", 10612 => "0010101100101000", 10613 => "1001111010111001", 10614 => "0100011111011000", 10615 => "0100000101111010", 10616 => "0010010100000100", 10617 => "0011100010011011", 10618 => "0100100100111001", 10619 => "0110011111101100", 10620 => "0111100101001010", 10621 => "0011001100001100", 10622 => "1111101010101000", 10623 => "0010110011101011", 10624 => "0010101011100100", 10625 => "0011011000100010", 10626 => "0011000110110001", 10627 => "1100110001011011", 10628 => "1001000101101011", 10629 => "1100101111000111", 10630 => "0010110000000101", 10631 => "0000110000010110", 10632 => "1110000101110101", 10633 => "0010111000010000", 10634 => "0000111011010011", 10635 => "1100010101110111", 10636 => "1101010011000001", 10637 => "0000110100001111", 10638 => "1010000110001000", 10639 => "1011011011000001", 10640 => "1010000110111100", 10641 => "1001111101011101", 10642 => "0001010111011000", 10643 => "0101011000001001", 10644 => "0110000110011111", 10645 => "0110011111001010", 10646 => "1110000011010010", 10647 => "0111101110111000", 10648 => "0011001111011011", 10649 => "1101000001011101", 10650 => "1000111101101010", 10651 => "1010000010101000", 10652 => "0000010001100001", 10653 => "0011000011101100", 10654 => "1000011010110001", 10655 => "0011101011110100", 10656 => "0100001101111011", 10657 => "1011011101011000", 10658 => "1010001000000100", 10659 => "1010101101100001", 10660 => "1011101011000010", 10661 => "0011111110010010", 10662 => "0110000010010111", 10663 => "1000100001000100", 10664 => "0001111001111011", 10665 => "1111010100111011", 10666 => "1010010110100100", 10667 => "1001101111101000", 10668 => "0001111000010100", 10669 => "1001010001001001", 10670 => "1101110001001101", 10671 => "1011001001101010", 10672 => "1100000110100101", 10673 => "0111111000011100", 10674 => "0100101011110001", 10675 => "1000010111111101", 10676 => "0000100000011011", 10677 => "0011101111001110", 10678 => "1100010000101000", 10679 => "0100110100010000", 10680 => "0011000011010100", 10681 => "1010101101011111", 10682 => "1010000111110100", 10683 => "1101110101101111", 10684 => "0101110101110101", 10685 => "1110110101010100", 10686 => "0011011011111110", 10687 => "0011101110111111", 10688 => "0111000001010001", 10689 => "1000111010010011", 10690 => "0011100101100011", 10691 => "0101011001010101", 10692 => "1111110101010001", 10693 => "1101110111011001", 10694 => "0101001111011011", 10695 => "1100110010011000", 10696 => "1001001010101110", 10697 => "0001010011010111", 10698 => "1011010011000111", 10699 => "1011100100111100", 10700 => "0011000010101111", 10701 => "0001010011011111", 10702 => "1111111001111010", 10703 => "0100001001100001", 10704 => "0111001111110110", 10705 => "0110001101111011", 10706 => "1100101100101001", 10707 => "0000010011110101", 10708 => "1100101100011010", 10709 => "0001010000101100", 10710 => "1000011111110101", 10711 => "1010110001010011", 10712 => "1001110011110111", 10713 => "1010111101011110", 10714 => "0001011010111101", 10715 => "1100001001111001", 10716 => "1011101000110101", 10717 => "1001000001100000", 10718 => "1110100111110111", 10719 => "1010110111100111", 10720 => "0100010010100011", 10721 => "0111111101110010", 10722 => "1100010100000011", 10723 => "0010100110000101", 10724 => "0111110001000100", 10725 => "0110001001101101", 10726 => "1000000001110110", 10727 => "1110111010010001", 10728 => "0110000100101110", 10729 => "0100100000110101", 10730 => "0010100101011100", 10731 => "1111101101100100", 10732 => "0000110011010110", 10733 => "0010000101100101", 10734 => "0110110000000010", 10735 => "0110111100101000", 10736 => "0101011111000110", 10737 => "0111001001110000", 10738 => "0001101010110001", 10739 => "1000111110001111", 10740 => "0011011001010110", 10741 => "1100111101001001", 10742 => "1010000011100111", 10743 => "1011101001010001", 10744 => "1100101101110100", 10745 => "0001001110110001", 10746 => "1101101100100000", 10747 => "0010100101001100", 10748 => "0100011111111011", 10749 => "0111000010100001", 10750 => "0111011010011000", 10751 => "1110101010001010", 10752 => "0010010100010010", 10753 => "1001100001011111", 10754 => "1000110011010110", 10755 => "0110001101110011", 10756 => "1100111101100011", 10757 => "0111100010011111", 10758 => "0100100101010000", 10759 => "1111111100011110", 10760 => "0000000100001110", 10761 => "0110001101100111", 10762 => "0000111100000110", 10763 => "1010001111100101", 10764 => "1011000100001011", 10765 => "1010011000101101", 10766 => "1111001011000101", 10767 => "1111011011011100", 10768 => "1100010100011010", 10769 => "0100110000010110", 10770 => "1001111100000110", 10771 => "0011001101111111", 10772 => "1110110011010110", 10773 => "1111111000100011", 10774 => "1101000101110011", 10775 => "0000100000010101", 10776 => "1011101000010010", 10777 => "0110101101100111", 10778 => "1101000010101111", 10779 => "1000010011000000", 10780 => "1001001000010001", 10781 => "1100011001100001", 10782 => "0001001010101101", 10783 => "0000011001111011", 10784 => "1111100010111111", 10785 => "1011011000001011", 10786 => "0001111001101101", 10787 => "1101000000011011", 10788 => "0101100001011001", 10789 => "1000110001010101", 10790 => "1101100110001000", 10791 => "1100111001000110", 10792 => "1111111101000101", 10793 => "1011101000100110", 10794 => "0100101000011000", 10795 => "0110000110011000", 10796 => "1100011011110010", 10797 => "0000100100111000", 10798 => "1111100100100010", 10799 => "1101110000111011", 10800 => "0011000100000110", 10801 => "1000100000110100", 10802 => "0101000000011010", 10803 => "1101001110011000", 10804 => "1000011111111010", 10805 => "0100101001011010", 10806 => "1011000001111111", 10807 => "0110111000110101", 10808 => "1011100001101100", 10809 => "0111111100000000", 10810 => "1001110111010110", 10811 => "0010100110100001", 10812 => "1011011001010110", 10813 => "1101000100111011", 10814 => "1011100001001011", 10815 => "0101011101001001", 10816 => "1110101100101101", 10817 => "0110110010000100", 10818 => "0100110011001110", 10819 => "1111110000110111", 10820 => "0100101011100101", 10821 => "0110101111010101", 10822 => "1011000101001100", 10823 => "1110100110000001", 10824 => "0110011100001110", 10825 => "1010101111101111", 10826 => "1001011110000101", 10827 => "0001110111001111", 10828 => "0010111100101100", 10829 => "1101111101111011", 10830 => "0010001000110111", 10831 => "1001000001110110", 10832 => "0010011111000111", 10833 => "1010010010000000", 10834 => "0011000000001001", 10835 => "1010111100011110", 10836 => "1011101101010000", 10837 => "0010011101010010", 10838 => "0010111100111110", 10839 => "0000111010001000", 10840 => "0110011100110011", 10841 => "1011101001111100", 10842 => "1111110001101110", 10843 => "0110101100111110", 10844 => "0100010110001100", 10845 => "1010001001001100", 10846 => "0011001111111111", 10847 => "1000110110100010", 10848 => "0000000010110001", 10849 => "1010101000110101", 10850 => "1111101110111100", 10851 => "1111001010110100", 10852 => "1101110011001001", 10853 => "0111000010101111", 10854 => "1100010001000111", 10855 => "0111100100011001", 10856 => "0110100110101100", 10857 => "0011001101001101", 10858 => "1100010111100100", 10859 => "1110010111010100", 10860 => "1110111111000011", 10861 => "1010001101111000", 10862 => "0101011110100000", 10863 => "1111100001101100", 10864 => "1001111000110010", 10865 => "1101001000011001", 10866 => "1101010101101111", 10867 => "1001001101101110", 10868 => "1101100010101110", 10869 => "0011110000100000", 10870 => "0001110111000011", 10871 => "1011101011110111", 10872 => "1001110100001110", 10873 => "1001100001100000", 10874 => "0111010100100010", 10875 => "0100010010111100", 10876 => "1100000000010010", 10877 => "0101111010110010", 10878 => "0010000000100010", 10879 => "0111010101100101", 10880 => "1100010010111100", 10881 => "1110100101010001", 10882 => "1111100001111001", 10883 => "0111101101110111", 10884 => "0101001001110101", 10885 => "1011011101000000", 10886 => "0000110111001111", 10887 => "0011010011100100", 10888 => "1010110110110111", 10889 => "1011010110100000", 10890 => "1100010000100000", 10891 => "0100100001111100", 10892 => "0101100101111011", 10893 => "1010100000001010", 10894 => "1010001000111101", 10895 => "1000111001010011", 10896 => "1001101010000111", 10897 => "0010111010110000", 10898 => "0101111001011111", 10899 => "1110111110000100", 10900 => "1101111100000110", 10901 => "0101000000101100", 10902 => "0001110000001111", 10903 => "1000010011001101", 10904 => "0111101010100001", 10905 => "1100110111010100", 10906 => "0010010000110011", 10907 => "1011100001101011", 10908 => "1110100000110011", 10909 => "0101110011110111", 10910 => "1110010110101011", 10911 => "1110011010011001", 10912 => "0110000000110111", 10913 => "1010111111001001", 10914 => "1010100001000111", 10915 => "1000010010101010", 10916 => "1101100001101110", 10917 => "0000001001011111", 10918 => "1101100010111111", 10919 => "1110010110100111", 10920 => "1001111000001011", 10921 => "0100110100001100", 10922 => "0001111100001110", 10923 => "0110010101010000", 10924 => "1000100010010110", 10925 => "0001101111100010", 10926 => "1011100101101001", 10927 => "0010010111000111", 10928 => "0001011111111011", 10929 => "1001010101011011", 10930 => "0110011011010111", 10931 => "0111011101011100", 10932 => "0001100001000100", 10933 => "1111110001110110", 10934 => "1000001010110101", 10935 => "0111000011001110", 10936 => "1001101100100001", 10937 => "1010101110111000", 10938 => "1000111010010011", 10939 => "0101110010011110", 10940 => "0010000101011101", 10941 => "1010110110101111", 10942 => "1111010011111011", 10943 => "0011101011100011", 10944 => "1100001110110000", 10945 => "1001001001110101", 10946 => "0101100011001001", 10947 => "0100011101000001", 10948 => "1001110001011101", 10949 => "0000001001101001", 10950 => "0101011000000000", 10951 => "0110010011101100", 10952 => "0101101001100010", 10953 => "0101001100011011", 10954 => "0001001111111100", 10955 => "1110001010011011", 10956 => "1110101001010000", 10957 => "1010000100111011", 10958 => "1000011111111011", 10959 => "1110100101001001", 10960 => "0110001000000110", 10961 => "1010011011101111", 10962 => "1001110000111110", 10963 => "0010011110100100", 10964 => "1000100010000001", 10965 => "0000100011101011", 10966 => "0100010100100010", 10967 => "0010001001110101", 10968 => "1101101011100001", 10969 => "0000110001010110", 10970 => "1000011000111001", 10971 => "0000111010111001", 10972 => "0110101010101100", 10973 => "0110000100000001", 10974 => "0111100110000001", 10975 => "0110100010110101", 10976 => "0111000001001101", 10977 => "0111111011110001", 10978 => "0100010111010010", 10979 => "1100111010111000", 10980 => "1001001100100100", 10981 => "0000010000010100", 10982 => "0010001110111110", 10983 => "0000101110000110", 10984 => "0111011100001101", 10985 => "1101101001111110", 10986 => "1110110100110011", 10987 => "0110011000100011", 10988 => "1110010100101010", 10989 => "1001010011011100", 10990 => "0111001100000010", 10991 => "1101111100100111", 10992 => "0000100000000110", 10993 => "1100111111100111", 10994 => "1100001101010100", 10995 => "0000110011000101", 10996 => "0111110101000010", 10997 => "0001110100111011", 10998 => "1010001000001101", 10999 => "0101101101010010", 11000 => "1101110110001000", 11001 => "0001000111101000", 11002 => "1110000001100010", 11003 => "1110010110101001", 11004 => "0111010000100110", 11005 => "0100110010001000", 11006 => "0011100011011001", 11007 => "1111101011110100", 11008 => "1111001011100010", 11009 => "1101000000000000", 11010 => "0001111111011100", 11011 => "1111000011011100", 11012 => "1001111011100111", 11013 => "0001011010111010", 11014 => "0011110100011001", 11015 => "1111100101011101", 11016 => "0000111110001101", 11017 => "1100110000100010", 11018 => "0001110001000100", 11019 => "0010000010011011", 11020 => "1110111011001011", 11021 => "1100010011000100", 11022 => "1010010110100010", 11023 => "0100010100001001", 11024 => "0011001110101110", 11025 => "1001011010011011", 11026 => "0100101010100111", 11027 => "0100110001011010", 11028 => "1101001011101100", 11029 => "1101000011111000", 11030 => "1101011111111100", 11031 => "1111000010100100", 11032 => "1010101101000000", 11033 => "0010110000100010", 11034 => "0011011111000011", 11035 => "0111011110100110", 11036 => "0000101101010011", 11037 => "1100010111101011", 11038 => "0001110101100010", 11039 => "0011101101100101", 11040 => "0000100001011001", 11041 => "1111001101100100", 11042 => "1100101111011000", 11043 => "1100000101111001", 11044 => "1100100111000000", 11045 => "0011100101000100", 11046 => "1000000101010010", 11047 => "1111010001111111", 11048 => "1100100100011011", 11049 => "1100010100000110", 11050 => "1101010010011100", 11051 => "0110000110001000", 11052 => "1000000110111101", 11053 => "1011000001110110", 11054 => "0100110000001011", 11055 => "1011111000010001", 11056 => "0011110110010011", 11057 => "0010010110010110", 11058 => "1111010100101001", 11059 => "1000101111110101", 11060 => "1101000101111000", 11061 => "0101101111001110", 11062 => "0011011101010110", 11063 => "1111000101000011", 11064 => "1001010011110110", 11065 => "0111010001001101", 11066 => "0100110000001110", 11067 => "1111100110110010", 11068 => "1101010001111111", 11069 => "0010100100110110", 11070 => "1100011010100001", 11071 => "1101100100110000", 11072 => "1111111101110111", 11073 => "0110010010100110", 11074 => "1000110001001100", 11075 => "0101101000010101", 11076 => "1100001001101011", 11077 => "1111100011011100", 11078 => "0000010100101001", 11079 => "0101111111111000", 11080 => "1011000111100010", 11081 => "0001001011000001", 11082 => "1100001100011001", 11083 => "1011110010001101", 11084 => "0100010101110100", 11085 => "1110001101011001", 11086 => "0011000010101010", 11087 => "0000111000011001", 11088 => "0000000010011110", 11089 => "1011110100010011", 11090 => "1110101001100101", 11091 => "0001010101001110", 11092 => "0110011010110010", 11093 => "0101101010110100", 11094 => "1000101101111000", 11095 => "0100100101010111", 11096 => "1010111110001010", 11097 => "0000011110111100", 11098 => "1001010100001110", 11099 => "1101100100001101", 11100 => "1001110010101101", 11101 => "1110010011100010", 11102 => "0100010101110010", 11103 => "0101000010010111", 11104 => "1011100000111010", 11105 => "1001101111110010", 11106 => "1111000010001101", 11107 => "1111110111001001", 11108 => "0000110111101111", 11109 => "0000101011001011", 11110 => "0110100000111110", 11111 => "1110100000000101", 11112 => "0001001111111111", 11113 => "0011101111011000", 11114 => "1110100111011000", 11115 => "1111110111011011", 11116 => "0000100010111001", 11117 => "1001100100111010", 11118 => "1000000100010110", 11119 => "1010000110000010", 11120 => "0101101000111001", 11121 => "0110100000000010", 11122 => "0010010110101001", 11123 => "1101111110000100", 11124 => "1001100100111111", 11125 => "0000111100011011", 11126 => "0000001011101010", 11127 => "1010011001011000", 11128 => "1000001100110001", 11129 => "0101011100100100", 11130 => "0010010011001111", 11131 => "0001110000001001", 11132 => "1000011111110001", 11133 => "0101111110001000", 11134 => "1100111001000101", 11135 => "1100101010010101", 11136 => "0110100000101101", 11137 => "1101110001101111", 11138 => "0010001100111100", 11139 => "0100001100110111", 11140 => "0001011000001001", 11141 => "1110010100111101", 11142 => "1101111101010110", 11143 => "0100110011010001", 11144 => "0101100100111000", 11145 => "1011110100110001", 11146 => "0111000110111101", 11147 => "1101010110011000", 11148 => "1011111011011111", 11149 => "1101010011100100", 11150 => "0010001011000011", 11151 => "0010001001000011", 11152 => "0111011110010101", 11153 => "1000001100110000", 11154 => "1000101110001110", 11155 => "1000110111001011", 11156 => "0110101000011110", 11157 => "0000001011110110", 11158 => "1000001000100000", 11159 => "0000111110001000", 11160 => "0011110011110110", 11161 => "0001001100110010", 11162 => "1101110000010011", 11163 => "0011011100010001", 11164 => "1000000001000111", 11165 => "1010010100101111", 11166 => "0101000101100100", 11167 => "0101011100001111", 11168 => "1111100011010001", 11169 => "0110101110000010", 11170 => "0010110111000111", 11171 => "0101000100111010", 11172 => "1100010100101101", 11173 => "0101011110111010", 11174 => "0110100011000111", 11175 => "0100010011001000", 11176 => "0000011011000011", 11177 => "0011100011111111", 11178 => "1111101110000101", 11179 => "0110101011001111", 11180 => "1010011011111110", 11181 => "1010011101001111", 11182 => "1010110110000000", 11183 => "0001100011110000", 11184 => "0000110010110110", 11185 => "1000001110010110", 11186 => "1010010000010000", 11187 => "0110001101101111", 11188 => "1000111001101100", 11189 => "1010001011111011", 11190 => "1110010111100111", 11191 => "1010101100111010", 11192 => "1010011111001100", 11193 => "0100101001110101", 11194 => "0001111100001110", 11195 => "0011111110101011", 11196 => "1010010011001100", 11197 => "1110000001010000", 11198 => "0000110010111001", 11199 => "1110000011000000", 11200 => "1010001100100001", 11201 => "0011001001001010", 11202 => "1111011010110010", 11203 => "1100011110010111", 11204 => "1010110100110100", 11205 => "1011100010011000", 11206 => "1000110001011000", 11207 => "1111010000001011", 11208 => "1010100001110010", 11209 => "1100110011001010", 11210 => "1000010011010111", 11211 => "0100000110110011", 11212 => "1100010111110000", 11213 => "0101101111111111", 11214 => "1000001110101001", 11215 => "1101101001001110", 11216 => "1000100101100010", 11217 => "0010011101000110", 11218 => "1001111111111110", 11219 => "0000110010011010", 11220 => "1100010110000111", 11221 => "0001110000111011", 11222 => "0010011110011101", 11223 => "0101111100111111", 11224 => "0011100101111110", 11225 => "1111100001000100", 11226 => "0100011101100010", 11227 => "1000010111110011", 11228 => "0011111010100001", 11229 => "0001010010011000", 11230 => "0111101010011001", 11231 => "1100010101111010", 11232 => "1000001100000101", 11233 => "1101011111000011", 11234 => "0111001100101000", 11235 => "0000001011111010", 11236 => "1010101000100011", 11237 => "1100100000010100", 11238 => "0111001011010001", 11239 => "1011001111101100", 11240 => "1100000110011110", 11241 => "1000111101110000", 11242 => "1100111110101011", 11243 => "0110010000011110", 11244 => "1010010111101101", 11245 => "1110000101100110", 11246 => "1111101011100011", 11247 => "0011010110101101", 11248 => "1100011011001010", 11249 => "1011000110100000", 11250 => "0100111011011110", 11251 => "1110011011000010", 11252 => "1100000000011100", 11253 => "1110011000110100", 11254 => "0001001110001001", 11255 => "0110001100010100", 11256 => "0100001101011000", 11257 => "0010110000100000", 11258 => "1011110111000010", 11259 => "1101110000101100", 11260 => "1010011000001011", 11261 => "1011010011101110", 11262 => "1010101001001110", 11263 => "0000001101111111", 11264 => "0101101101000101", 11265 => "0100011000101111", 11266 => "0011011010110110", 11267 => "1000001111111001", 11268 => "0111011101111110", 11269 => "1000000100011100", 11270 => "0101100001110010", 11271 => "1110101010100110", 11272 => "1111110010001011", 11273 => "0010010010110110", 11274 => "0010110001010100", 11275 => "0001110111001001", 11276 => "0101000010011110", 11277 => "0010100100000011", 11278 => "0100110001001010", 11279 => "1001000110100110", 11280 => "1011000001100010", 11281 => "1110001101001010", 11282 => "1111100001011001", 11283 => "0110111000011010", 11284 => "1000101100011111", 11285 => "1100110000100111", 11286 => "1100101011111101", 11287 => "1101001001110000", 11288 => "0110101000111000", 11289 => "1000100110110011", 11290 => "1011101011110000", 11291 => "1101101110011100", 11292 => "0010100110011010", 11293 => "0001100111000100", 11294 => "0100100111010001", 11295 => "1000111001111010", 11296 => "1101101001100011", 11297 => "0110110010010001", 11298 => "0100100010010001", 11299 => "0011011011001111", 11300 => "0111010100000100", 11301 => "0001101001001100", 11302 => "0001110000101010", 11303 => "0011001100101001", 11304 => "0100000001001000", 11305 => "0110100000101000", 11306 => "1000101110101101", 11307 => "0111011010111011", 11308 => "1110100010111111", 11309 => "0100001111101010", 11310 => "0010000001110010", 11311 => "1101010110001000", 11312 => "1001011111001000", 11313 => "1010110100010111", 11314 => "1110001011010111", 11315 => "0110010110100111", 11316 => "0011111100011111", 11317 => "1110010111010010", 11318 => "1110101110000011", 11319 => "1000100011011010", 11320 => "0001010001000010", 11321 => "0111100010101100", 11322 => "0011001011110001", 11323 => "0100000010010001", 11324 => "1001101110010101", 11325 => "1111011101111110", 11326 => "0111000100011010", 11327 => "1110000010001100", 11328 => "1100111101100111", 11329 => "0011010011000011", 11330 => "0110110101110011", 11331 => "1111001101110000", 11332 => "0101111110101111", 11333 => "0010101110010011", 11334 => "1001111010110101", 11335 => "0001010110110110", 11336 => "1111111000000010", 11337 => "1011001101100111", 11338 => "1111011110101000", 11339 => "0100101101101010", 11340 => "0011111111110000", 11341 => "0110011010011111", 11342 => "0110110001111010", 11343 => "1100011000010111", 11344 => "0100011000110011", 11345 => "1100100100010001", 11346 => "0101011010100100", 11347 => "0100011111100001", 11348 => "1000010111101011", 11349 => "1100111111101111", 11350 => "0000101110110001", 11351 => "0010010111100100", 11352 => "1110101110101000", 11353 => "0101110011111011", 11354 => "1010110111000001", 11355 => "0011101010111000", 11356 => "0101110100111101", 11357 => "0001100100011100", 11358 => "1010111000000011", 11359 => "1010010000101110", 11360 => "1110100001110000", 11361 => "0100000010100110", 11362 => "0101001000111101", 11363 => "0000011010001000", 11364 => "0011000110000111", 11365 => "0000111101111100", 11366 => "0011111101001000", 11367 => "1111101001101100", 11368 => "1111001111011110", 11369 => "0101100010100010", 11370 => "1100101000100101", 11371 => "0100011011000011", 11372 => "0111101101110010", 11373 => "1010000101011011", 11374 => "0000110001100101", 11375 => "1110100110100100", 11376 => "1010001010011101", 11377 => "1100000001101011", 11378 => "0001011101100111", 11379 => "0101111111011001", 11380 => "1110100010101001", 11381 => "1001111101100001", 11382 => "0000100001000001", 11383 => "1011111010010001", 11384 => "1110101000111001", 11385 => "1110110110101011", 11386 => "1100110100111010", 11387 => "1011101100101011", 11388 => "0001010101111100", 11389 => "0101111101101100", 11390 => "0110000111001011", 11391 => "0110111110011110", 11392 => "1011010101100010", 11393 => "1110110111111010", 11394 => "1111000101010101", 11395 => "1010010110001111", 11396 => "1001111011101101", 11397 => "0010001011101100", 11398 => "1000110011110101", 11399 => "1001011111110100", 11400 => "1110000001011101", 11401 => "1110111001110100", 11402 => "0010111001011111", 11403 => "0010000010111011", 11404 => "1010100001010111", 11405 => "1101000011110100", 11406 => "1110000010110100", 11407 => "1111011011010001", 11408 => "1011110101111010", 11409 => "1110111010110001", 11410 => "0111010100100110", 11411 => "0000000100011000", 11412 => "1110001001100111", 11413 => "1101001110110000", 11414 => "1000111011101101", 11415 => "0110111111010101", 11416 => "0101000010001100", 11417 => "1101011001101010", 11418 => "0101101110010101", 11419 => "0110001110010011", 11420 => "0000011100110110", 11421 => "1111000100100110", 11422 => "0000000101000100", 11423 => "0010100111011111", 11424 => "1111000111101110", 11425 => "0000001010101001", 11426 => "0011010111011010", 11427 => "1010111000001001", 11428 => "1111001111110001", 11429 => "1000111000101101", 11430 => "1110110111101111", 11431 => "0100011000110011", 11432 => "1101000010001000", 11433 => "1001010111000000", 11434 => "0000010001100100", 11435 => "0100011100101000", 11436 => "1011010110010100", 11437 => "1110101110110110", 11438 => "1111111010010111", 11439 => "0000110110011100", 11440 => "1100111111111011", 11441 => "1000010101010001", 11442 => "1101100011100010", 11443 => "0000110100111111", 11444 => "1110110001100010", 11445 => "0000100010000010", 11446 => "0011011001111110", 11447 => "0110101110000000", 11448 => "1110100101001101", 11449 => "1110100100010110", 11450 => "0110011011101111", 11451 => "1101110000001010", 11452 => "0001000111010110", 11453 => "1001110011101101", 11454 => "0010011011011011", 11455 => "1011010010100001", 11456 => "1110111011010101", 11457 => "1110100000011110", 11458 => "0101001000010001", 11459 => "1110001011101001", 11460 => "0010000010110011", 11461 => "1000001000010110", 11462 => "0100000001101110", 11463 => "0010111100001001", 11464 => "1010001110101101", 11465 => "1000010111110011", 11466 => "0000101011011110", 11467 => "0110011010000101", 11468 => "0101000111110111", 11469 => "0010100010000101", 11470 => "0100000111111000", 11471 => "0100110011101000", 11472 => "0000100100110001", 11473 => "1010011110110010", 11474 => "1111110000011100", 11475 => "0001010001011011", 11476 => "1001010100110001", 11477 => "1000001100001111", 11478 => "1110110111101001", 11479 => "0110000110010100", 11480 => "0000100110111111", 11481 => "1111011101110101", 11482 => "0011100101110000", 11483 => "1010010100100011", 11484 => "0000000111000100", 11485 => "0101110010111001", 11486 => "0010100101000100", 11487 => "0000000111111011", 11488 => "1100010111111001", 11489 => "1001010000101010", 11490 => "0000000101100001", 11491 => "1110111101101011", 11492 => "0100111000011111", 11493 => "1010100000001110", 11494 => "0011010010100101", 11495 => "0100000110001111", 11496 => "1011000010000011", 11497 => "0011101101111111", 11498 => "1001111010101001", 11499 => "1110110001100010", 11500 => "1000001101110001", 11501 => "0111001000001111", 11502 => "1011110100000101", 11503 => "0111100100110000", 11504 => "0001010101101011", 11505 => "0000101001100101", 11506 => "0000100010111111", 11507 => "0100100100001011", 11508 => "0110000101101100", 11509 => "1101111101100101", 11510 => "1001101110110100", 11511 => "0011100000111111", 11512 => "0100111110100011", 11513 => "1100111100000110", 11514 => "1010000100000100", 11515 => "1111000010010010", 11516 => "1110111001010001", 11517 => "0100110000111011", 11518 => "1011000011101000", 11519 => "1111100010000100", 11520 => "0110000100110000", 11521 => "1000010111010110", 11522 => "1001010010000110", 11523 => "0100100001111111", 11524 => "1111011110010100", 11525 => "0011011010001111", 11526 => "0000010010011010", 11527 => "1101110111001101", 11528 => "1110000110100000", 11529 => "1110000001101100", 11530 => "0011100100100011", 11531 => "1011111001000000", 11532 => "1011111110111011", 11533 => "0111111010011001", 11534 => "1101001011010011", 11535 => "1011110100000000", 11536 => "1011011110101100", 11537 => "0000111111011101", 11538 => "0111101101100101", 11539 => "1011110110000001", 11540 => "0100101100110100", 11541 => "1001011000011111", 11542 => "0000011001010011", 11543 => "0000000010110011", 11544 => "0010011100111111", 11545 => "1000110000011101", 11546 => "0000111010100100", 11547 => "1000001100000101", 11548 => "0111010110100011", 11549 => "1010101100000000", 11550 => "0001000010100010", 11551 => "0110111001011101", 11552 => "0010001110101011", 11553 => "1100001110101011", 11554 => "0010001111010000", 11555 => "0001011100110111", 11556 => "0010010001100011", 11557 => "0011001111100001", 11558 => "1101000010011110", 11559 => "0100000010110100", 11560 => "1111101111001111", 11561 => "1000001100000100", 11562 => "1100110110001110", 11563 => "1100111101010000", 11564 => "0101010011010010", 11565 => "0000000111100111", 11566 => "0001101100101011", 11567 => "0011000011001110", 11568 => "1110010100001100", 11569 => "0011001000101100", 11570 => "0010110111101110", 11571 => "1010110110010000", 11572 => "0101001000111011", 11573 => "0011100101000011", 11574 => "1001011011111001", 11575 => "0000000101010010", 11576 => "1101010100111010", 11577 => "1011111010111010", 11578 => "1000000000010011", 11579 => "1100010001010111", 11580 => "0111001101110100", 11581 => "0111011011000110", 11582 => "0110011111111110", 11583 => "0000001011011000", 11584 => "0001000101101011", 11585 => "1101001100011110", 11586 => "0011110110101011", 11587 => "1000011000110011", 11588 => "1111111011001110", 11589 => "1110011001111111", 11590 => "1110001010001010", 11591 => "1000100011000111", 11592 => "1100101101001100", 11593 => "1001101111000001", 11594 => "1011101010010101", 11595 => "0101110000101111", 11596 => "1100111011111001", 11597 => "0000001101011001", 11598 => "1011011010101111", 11599 => "0011101001001111", 11600 => "0011100111010110", 11601 => "1111101010000101", 11602 => "0011110000001000", 11603 => "1000110010111011", 11604 => "0000001100001010", 11605 => "1010101000010111", 11606 => "1110011110110100", 11607 => "0110010101100011", 11608 => "1000001111111000", 11609 => "0000111111100110", 11610 => "0110000100010101", 11611 => "0110010011011100", 11612 => "1001011000001000", 11613 => "1111000100101011", 11614 => "1111100010010111", 11615 => "0100010110011011", 11616 => "0001101000000010", 11617 => "1110010001010100", 11618 => "0100111001110110", 11619 => "0100000101001110", 11620 => "1010100001101111", 11621 => "1111101100101110", 11622 => "0101110110111100", 11623 => "1000110100110110", 11624 => "0010101010000001", 11625 => "0011101110101100", 11626 => "1000010001000111", 11627 => "0000111111000000", 11628 => "0000010101000010", 11629 => "0011010100110010", 11630 => "1001110011111000", 11631 => "0010011100010000", 11632 => "1100000110101011", 11633 => "1101101100001001", 11634 => "0110111001001100", 11635 => "1010110100000110", 11636 => "1100011011000101", 11637 => "1010111010110111", 11638 => "1010100010100010", 11639 => "0011110000101110", 11640 => "1110111111011001", 11641 => "1011111010111010", 11642 => "1010001100001001", 11643 => "1000101000001101", 11644 => "1000110110000011", 11645 => "0101001101010010", 11646 => "0100100011110100", 11647 => "0101111110000010", 11648 => "1000001001010011", 11649 => "1001111010000000", 11650 => "1001100011100000", 11651 => "0010100000110100", 11652 => "0100000010101011", 11653 => "0110001011010000", 11654 => "1100001001110100", 11655 => "1011110110000111", 11656 => "1111111001011111", 11657 => "1011110000010011", 11658 => "0001100101111011", 11659 => "0110100100000110", 11660 => "0111000001001110", 11661 => "0010100101000000", 11662 => "0010010000001010", 11663 => "1111010010011100", 11664 => "1010000101110110", 11665 => "0101110111010100", 11666 => "0111101110100000", 11667 => "0110111110101111", 11668 => "0101100111010000", 11669 => "1100001111100001", 11670 => "0010000011000101", 11671 => "1010111000111101", 11672 => "0111101000010000", 11673 => "1001011011010010", 11674 => "0100001100100000", 11675 => "1000101011100001", 11676 => "1011100011111011", 11677 => "1110001001101100", 11678 => "0111101101011010", 11679 => "0000001101001011", 11680 => "0101000111010011", 11681 => "0011110000100000", 11682 => "1001110000110000", 11683 => "1011000111010011", 11684 => "1010101000111101", 11685 => "1100011111100001", 11686 => "0000101100110100", 11687 => "1010010110101000", 11688 => "1110000011011110", 11689 => "0101001111111010", 11690 => "0010011001101111", 11691 => "0111011010001101", 11692 => "1011101111011000", 11693 => "0111111100000001", 11694 => "0111100010101101", 11695 => "0010101001101100", 11696 => "0011101010101000", 11697 => "1111101101001101", 11698 => "1100001100101001", 11699 => "1000100010101000", 11700 => "1010111010010111", 11701 => "1010111100111001", 11702 => "0111111010010011", 11703 => "0010110100101101", 11704 => "0000001010111111", 11705 => "0111110000000001", 11706 => "1100101111000110", 11707 => "1000011000011111", 11708 => "1111000111101110", 11709 => "0011101001100011", 11710 => "1111111010110110", 11711 => "1011011100011000", 11712 => "0001010000100010", 11713 => "0010111110011000", 11714 => "1011100101001000", 11715 => "1111000000111001", 11716 => "1101110001011100", 11717 => "1000110111100100", 11718 => "0111100010101000", 11719 => "0000000100110000", 11720 => "1001111100110101", 11721 => "1000010001001100", 11722 => "1100110110100000", 11723 => "1111101100010111", 11724 => "0110110001001001", 11725 => "1001111100110001", 11726 => "1011001000010110", 11727 => "0011110000001110", 11728 => "1110110110011110", 11729 => "0111100101011111", 11730 => "0000101000110110", 11731 => "1001001110110000", 11732 => "1010101101000110", 11733 => "0000101111000011", 11734 => "1010110000101011", 11735 => "0110101011011101", 11736 => "1111010101110000", 11737 => "1010001010101100", 11738 => "1100001010010100", 11739 => "0110010111001101", 11740 => "0010000011100110", 11741 => "0111001010001001", 11742 => "1110101001111000", 11743 => "1110011010010000", 11744 => "1111111101111111", 11745 => "1101100010010011", 11746 => "0001011110101010", 11747 => "1000101010011111", 11748 => "0010000000011000", 11749 => "1111000000010010", 11750 => "1110010111101011", 11751 => "1110110010001101", 11752 => "1011101101101011", 11753 => "1111000001001000", 11754 => "1101001100000010", 11755 => "0001111011111111", 11756 => "0100100101110100", 11757 => "0110010111010011", 11758 => "1011000110101110", 11759 => "1101001101101000", 11760 => "0001110000110001", 11761 => "0100011111110100", 11762 => "0001011001110000", 11763 => "0001000000000010", 11764 => "1011000010001101", 11765 => "0100111000011101", 11766 => "0111111011110111", 11767 => "0010010011000111", 11768 => "1001000110111010", 11769 => "0000000101010011", 11770 => "0111001100101011", 11771 => "1111000100101101", 11772 => "0000111000100001", 11773 => "0110110000100101", 11774 => "0000001110010111", 11775 => "0010001000000001", 11776 => "0101110110110011", 11777 => "0100011001111101", 11778 => "1101001010010110", 11779 => "1110100010000101", 11780 => "0101101010010011", 11781 => "0000111101010100", 11782 => "1010001100010000", 11783 => "0111101110001001", 11784 => "0110101100110100", 11785 => "0000001101011101", 11786 => "0001010101101101", 11787 => "0100001011100101", 11788 => "1001100010111001", 11789 => "0001011011100101", 11790 => "0110001100011101", 11791 => "0110010001110100", 11792 => "0000100101011001", 11793 => "1000001111100010", 11794 => "0010010000111101", 11795 => "1001010100011000", 11796 => "1110000010010100", 11797 => "0111010010101010", 11798 => "1011101000011101", 11799 => "1011010101000001", 11800 => "0100101011000100", 11801 => "0111010000011101", 11802 => "1010101011110111", 11803 => "1111000111101001", 11804 => "1111100100100010", 11805 => "0110000111100000", 11806 => "0010110111100010", 11807 => "1100111001101111", 11808 => "1111110000100111", 11809 => "1011111001110101", 11810 => "1010110101111011", 11811 => "0110011111110111", 11812 => "0010111010001010", 11813 => "0101010110011011", 11814 => "1111110111010001", 11815 => "1011001110100011", 11816 => "1111101110000100", 11817 => "1111101001100011", 11818 => "0101011101001010", 11819 => "0000100110110110", 11820 => "1001010010000000", 11821 => "1111001111010010", 11822 => "1001000011110000", 11823 => "0100010110011101", 11824 => "0110110100011000", 11825 => "0100111101000101", 11826 => "1011110100011011", 11827 => "1100101101111101", 11828 => "0011010110100110", 11829 => "1010001101010000", 11830 => "1100000010000110", 11831 => "1011001101110111", 11832 => "1110010110010011", 11833 => "1111001111000001", 11834 => "0001011010011011", 11835 => "0101000110011001", 11836 => "1010010111010100", 11837 => "0010110111111110", 11838 => "0000010101110101", 11839 => "0101101110011011", 11840 => "0011101011101110", 11841 => "0110110010110111", 11842 => "1011000010100010", 11843 => "0001001001101011", 11844 => "0101001011100101", 11845 => "0100000001001010", 11846 => "1001000011100110", 11847 => "0110011101100110", 11848 => "0010001101011011", 11849 => "1001101110110000", 11850 => "1111001010100010", 11851 => "0111101100101000", 11852 => "0010011001101100", 11853 => "0111011000011010", 11854 => "1010000111001111", 11855 => "0011010000010100", 11856 => "0001011011011110", 11857 => "0001100101010110", 11858 => "0111010010011000", 11859 => "0110110001110001", 11860 => "0101001010110101", 11861 => "1010110111100110", 11862 => "0100110101011111", 11863 => "1101010100100010", 11864 => "1100011110000001", 11865 => "0101001010101011", 11866 => "1000100111111110", 11867 => "0110100100100000", 11868 => "1000101001101110", 11869 => "0100010100110000", 11870 => "0011100001110111", 11871 => "1000011000010000", 11872 => "0100101101110010", 11873 => "0110101101001001", 11874 => "1011001011101011", 11875 => "1010100111001000", 11876 => "0010101100111101", 11877 => "0010101100101101", 11878 => "1111110010010110", 11879 => "0111010000111111", 11880 => "1100110000011110", 11881 => "0010100011000010", 11882 => "0101110010000100", 11883 => "1001110011001110", 11884 => "0010101111100001", 11885 => "0010001100111010", 11886 => "0101111010000101", 11887 => "0100001011001111", 11888 => "0011000110100110", 11889 => "1010101110010111", 11890 => "1111001011100010", 11891 => "1010001101010100", 11892 => "0110011010100110", 11893 => "1111011101100110", 11894 => "1101111001110000", 11895 => "0100101000101101", 11896 => "1100001110001100", 11897 => "0000111001001011", 11898 => "1001111100010110", 11899 => "1010001000101001", 11900 => "1010000011010111", 11901 => "1000011110000010", 11902 => "1010001110110111", 11903 => "0001001111001011", 11904 => "1100010101001100", 11905 => "0101101010011110", 11906 => "0001000010010111", 11907 => "0011001111001001", 11908 => "0100000001010111", 11909 => "1101010010110101", 11910 => "0101100001011100", 11911 => "0110000001010001", 11912 => "0001101110000100", 11913 => "1110111111011110", 11914 => "1010010010000011", 11915 => "1110010101000010", 11916 => "1110001001010001", 11917 => "1010000010011101", 11918 => "0000001110111101", 11919 => "1001001010000101", 11920 => "1101011001111111", 11921 => "1011010101011000", 11922 => "0101000101101010", 11923 => "1100110000110111", 11924 => "1001110011111100", 11925 => "1111111011100000", 11926 => "0011000011110100", 11927 => "0011000101110100", 11928 => "0111110011110111", 11929 => "0111011100110011", 11930 => "0001110001011101", 11931 => "0001100101100101", 11932 => "1010000010100011", 11933 => "0101101010111000", 11934 => "1111101000001111", 11935 => "1111011100110000", 11936 => "1101010011111011", 11937 => "1101100010110110", 11938 => "0100001110111010", 11939 => "0110000100101011", 11940 => "0010011100011101", 11941 => "1101100011001110", 11942 => "0010101010011000", 11943 => "0100100010011010", 11944 => "1010100111000011", 11945 => "0001111010010001", 11946 => "1011000010101001", 11947 => "0001110111111010", 11948 => "1100010011101010", 11949 => "1000110000011001", 11950 => "0100101111101111", 11951 => "1001110110011000", 11952 => "1110010110000100", 11953 => "0110111111111001", 11954 => "0011001101010101", 11955 => "0100010011111000", 11956 => "1111100110011001", 11957 => "0011110000101101", 11958 => "1100101001100100", 11959 => "1011010010101111", 11960 => "1011001001100010", 11961 => "0001110011101100", 11962 => "0101111100000000", 11963 => "1111001000110101", 11964 => "1101011010101111", 11965 => "1101110000011100", 11966 => "0011100001001110", 11967 => "0000001100010100", 11968 => "1111011101101100", 11969 => "1101001001000001", 11970 => "0000001001011001", 11971 => "1101110010111100", 11972 => "1001000111110111", 11973 => "0010000011110011", 11974 => "1011101110110011", 11975 => "1110010100010110", 11976 => "1011111010000110", 11977 => "1000000110101010", 11978 => "1000101110110001", 11979 => "0101111100001001", 11980 => "1010011100010010", 11981 => "1110000010010000", 11982 => "1101000100011001", 11983 => "1101100011101001", 11984 => "1000010011001111", 11985 => "1010101001000011", 11986 => "1011100111110100", 11987 => "0010101100001010", 11988 => "1100010001101101", 11989 => "1100101000110111", 11990 => "0000010110010110", 11991 => "0101000001100111", 11992 => "1100100001001110", 11993 => "1010010001111111", 11994 => "0100110111010111", 11995 => "1101011110011010", 11996 => "0101011100100010", 11997 => "0010100100111101", 11998 => "1001001111010011", 11999 => "1111111110101001", 12000 => "0110101110101100", 12001 => "1010000111100010", 12002 => "1101110000101011", 12003 => "1001010101101010", 12004 => "1111011011101010", 12005 => "1111110001101100", 12006 => "0011101101000110", 12007 => "1000111101101101", 12008 => "1000011100111001", 12009 => "1111001000000100", 12010 => "1000100000011011", 12011 => "0111111001100111", 12012 => "0000011001111110", 12013 => "1101010000001001", 12014 => "1001110011101000", 12015 => "0001011110100101", 12016 => "1100111110000101", 12017 => "1010111100010000", 12018 => "0110000110110111", 12019 => "1000110111000010", 12020 => "1011110000100010", 12021 => "1000110110110110", 12022 => "0110011010101010", 12023 => "1011011011011101", 12024 => "0101110100101100", 12025 => "1001110100110011", 12026 => "1110000110011010", 12027 => "0001100111000111", 12028 => "0001110011110111", 12029 => "0111110100110111", 12030 => "1000100100001001", 12031 => "0101011111011100", 12032 => "0010101001111001", 12033 => "0010000110010011", 12034 => "0001100000100111", 12035 => "1001001000110000", 12036 => "0100111011001100", 12037 => "0001011000011100", 12038 => "0110010011101111", 12039 => "0100111001111010", 12040 => "0000010000000011", 12041 => "1010101011001001", 12042 => "0011010010000010", 12043 => "1010100001010101", 12044 => "1111111001111110", 12045 => "0110010001001000", 12046 => "1011110111000010", 12047 => "0000111111111010", 12048 => "1110111110010001", 12049 => "0001111101001110", 12050 => "1001100010011010", 12051 => "0001011010010111", 12052 => "1011001100101001", 12053 => "1011011110001100", 12054 => "1011100101010001", 12055 => "1111001010000011", 12056 => "1110011101110111", 12057 => "0110011000001001", 12058 => "1110101011001001", 12059 => "0110110101111110", 12060 => "0111100111010000", 12061 => "1101000001100010", 12062 => "1110110000000110", 12063 => "0110101001111011", 12064 => "1010100010001001", 12065 => "1001000000111000", 12066 => "0001100010101001", 12067 => "0010101110101111", 12068 => "1110110110000101", 12069 => "1000101101101010", 12070 => "0110101010011100", 12071 => "0111111100001110", 12072 => "1110110111100111", 12073 => "0110100110101001", 12074 => "1111010111101100", 12075 => "0110100010100101", 12076 => "0010010001001010", 12077 => "1011101010000010", 12078 => "0100110000111101", 12079 => "1110011000011101", 12080 => "1110111000010100", 12081 => "1100100001100110", 12082 => "0111111011101000", 12083 => "0100111101010000", 12084 => "1010000011110011", 12085 => "1000000010101101", 12086 => "1100110111100010", 12087 => "0100110010000111", 12088 => "1000100000100111", 12089 => "1110011001011001", 12090 => "0100001111001001", 12091 => "1101011010111010", 12092 => "1100100001011010", 12093 => "1110001001001101", 12094 => "1110111100010001", 12095 => "1000111100001101", 12096 => "1010101001101011", 12097 => "0110111110000011", 12098 => "1111110101110110", 12099 => "0010010001101110", 12100 => "1011011100101110", 12101 => "0011010100101100", 12102 => "0111000111011000", 12103 => "1011010000101100", 12104 => "0101001111110110", 12105 => "1011101111000110", 12106 => "1011110111110100", 12107 => "0000100011010010", 12108 => "0000101010001111", 12109 => "1011001001000010", 12110 => "1011111101011011", 12111 => "0010110001000101", 12112 => "0110111101100100", 12113 => "1101101110011010", 12114 => "0010001000111000", 12115 => "0110110010100100", 12116 => "1001010011010100", 12117 => "1010110101000001", 12118 => "1110010100100010", 12119 => "1001000010010100", 12120 => "0111000010100100", 12121 => "0101010110111011", 12122 => "1110110111100000", 12123 => "1010001110000000", 12124 => "1100010011111110", 12125 => "0010000111010010", 12126 => "0010010010010101", 12127 => "1110010111001000", 12128 => "0011011001100101", 12129 => "1010111111110001", 12130 => "0000110110110100", 12131 => "0111101101101100", 12132 => "1011101111101001", 12133 => "1001101101001011", 12134 => "0101110100000000", 12135 => "0010011001000110", 12136 => "1011010001111000", 12137 => "1100000110111111", 12138 => "1101110001010100", 12139 => "0110010000101001", 12140 => "1010010001000000", 12141 => "1100001101010100", 12142 => "1011000000101001", 12143 => "0001001001001001", 12144 => "1001101010110001", 12145 => "1111011001100011", 12146 => "1100110001010001", 12147 => "1001111111010001", 12148 => "1000100011101100", 12149 => "1110010100100000", 12150 => "1000000110010110", 12151 => "0101000100010001", 12152 => "0011011000111000", 12153 => "0011111101000000", 12154 => "1111110100000001", 12155 => "1000100101011101", 12156 => "1110111110010101", 12157 => "0101001111100110", 12158 => "0011100100111001", 12159 => "1111111001010011", 12160 => "1011010010110101", 12161 => "0100000011000110", 12162 => "0001011111001011", 12163 => "0101100110011100", 12164 => "0100110000010100", 12165 => "1111101100011101", 12166 => "0000001100101100", 12167 => "1011101100100101", 12168 => "0010100110010011", 12169 => "0101001001111101", 12170 => "1011111011011011", 12171 => "1101001000101000", 12172 => "1100101101011001", 12173 => "0000100010101001", 12174 => "1010001101110001", 12175 => "1101010010010101", 12176 => "0110010001101000", 12177 => "1101111110000111", 12178 => "1010100111010101", 12179 => "1001011111010110", 12180 => "1110110001011101", 12181 => "0110101100111001", 12182 => "1000011111110001", 12183 => "1110001011010111", 12184 => "0010111101010000", 12185 => "1001000011001001", 12186 => "0110000010000110", 12187 => "0110110110001011", 12188 => "1101101011111111", 12189 => "0011101110110001", 12190 => "0000110100110001", 12191 => "1011001110010110", 12192 => "1100100101100101", 12193 => "0000111111000111", 12194 => "1101010010001101", 12195 => "0000010101011111", 12196 => "0001000001010100", 12197 => "1000111001011010", 12198 => "0000110011100010", 12199 => "0101010110001001", 12200 => "1111000000111011", 12201 => "1101011110101110", 12202 => "0010101111100011", 12203 => "1111111101101111", 12204 => "0011001001100001", 12205 => "1010101100100111", 12206 => "1100011011111010", 12207 => "1010010100100100", 12208 => "1011101011010011", 12209 => "1101101000101000", 12210 => "0000110110110100", 12211 => "0110000100110000", 12212 => "1001000001001010", 12213 => "1000110100011000", 12214 => "0001110110000000", 12215 => "0111000110011110", 12216 => "1111011001100100", 12217 => "0110110001111101", 12218 => "0111010010111010", 12219 => "0011110110001001", 12220 => "1010010110100010", 12221 => "0101000011111100", 12222 => "0110100110010010", 12223 => "0010111100011110", 12224 => "1111110100100010", 12225 => "1011010011001100", 12226 => "1010011010011010", 12227 => "1000011111110011", 12228 => "1111111011110001", 12229 => "0011001000000010", 12230 => "0100110010010000", 12231 => "0100110000001100", 12232 => "0110001010010000", 12233 => "0110100001001001", 12234 => "0101011101111101", 12235 => "0010110000111101", 12236 => "0011010111011100", 12237 => "0101111101010100", 12238 => "1101111011010001", 12239 => "1001011101111111", 12240 => "0011101100011101", 12241 => "1100100100101111", 12242 => "0110100100100010", 12243 => "0010000011111110", 12244 => "0110010010110110", 12245 => "0001111111000111", 12246 => "1100110010101000", 12247 => "1000001010101111", 12248 => "0110010110001101", 12249 => "1100101010010000", 12250 => "0111110010011011", 12251 => "1010100100110001", 12252 => "0100010010001111", 12253 => "0100000010111000", 12254 => "1111111000110100", 12255 => "1111100101100101", 12256 => "1011100011011101", 12257 => "0000111111011110", 12258 => "1111000011001111", 12259 => "1100011011110011", 12260 => "0100001100100010", 12261 => "1111001100101001", 12262 => "1101011001011110", 12263 => "0010100000010111", 12264 => "0111111111011011", 12265 => "1000100000011111", 12266 => "1011000001110001", 12267 => "1011010011011011", 12268 => "0000110110000010", 12269 => "0100101111011000", 12270 => "1101010001010111", 12271 => "0001111100010100", 12272 => "0101111011010110", 12273 => "1111001100101110", 12274 => "0011111100111101", 12275 => "1000011011101111", 12276 => "0100001110110010", 12277 => "1111111000101010", 12278 => "0110111011110100", 12279 => "1111101011111111", 12280 => "0101110001101000", 12281 => "0100110001011001", 12282 => "1001000001011101", 12283 => "0011111011110110", 12284 => "0100110111011101", 12285 => "1101010001111000", 12286 => "0110011110001011", 12287 => "1110110110100110", 12288 => "1000000011010000", 12289 => "0010001100000011", 12290 => "1000011000110001", 12291 => "1110100111111100", 12292 => "0001010001100011", 12293 => "0110011001011100", 12294 => "0100010111000111", 12295 => "0111001010000000", 12296 => "1110111101110000", 12297 => "1011110011011101", 12298 => "0011111010011010", 12299 => "1000001110100001", 12300 => "1011001111100100", 12301 => "1101110001001010", 12302 => "0100010001111111", 12303 => "0000101111010001", 12304 => "1111111101010001", 12305 => "0011100111001101", 12306 => "0100011000101010", 12307 => "1101000111100111", 12308 => "1111111011110100", 12309 => "1111011001001111", 12310 => "1110100000011100", 12311 => "1110011100010100", 12312 => "0110010110101011", 12313 => "0111011011111110", 12314 => "0011010010100001", 12315 => "1011111101010110", 12316 => "0100011001011011", 12317 => "1011011101101011", 12318 => "0000111100000110", 12319 => "0100010011000010", 12320 => "0011100110110101", 12321 => "1000010110101100", 12322 => "0011010110101001", 12323 => "1110001011100110", 12324 => "1101101010100011", 12325 => "0101001001101111", 12326 => "0110001000000010", 12327 => "0100011011111010", 12328 => "0000011001001011", 12329 => "0101010001110000", 12330 => "1111001001000000", 12331 => "0001011001100100", 12332 => "1111110100110100", 12333 => "1000010101001110", 12334 => "0110000100000100", 12335 => "0001001111110101", 12336 => "1000111101101011", 12337 => "0100000110011000", 12338 => "1111101110111100", 12339 => "1000100001011101", 12340 => "1000011000100001", 12341 => "0111100001001100", 12342 => "0011101100101010", 12343 => "1100001011011101", 12344 => "1011011010110100", 12345 => "0100010110111110", 12346 => "0111110110011110", 12347 => "1011100100111110", 12348 => "0011000110110101", 12349 => "1101110010011000", 12350 => "0001001111010011", 12351 => "0000100100101110", 12352 => "1001000010001011", 12353 => "0110001010000110", 12354 => "0101011000001111", 12355 => "1111011000111100", 12356 => "0001000011111000", 12357 => "0101011000101100", 12358 => "0101100011001010", 12359 => "1111100101011100", 12360 => "0101100010000011", 12361 => "0011010100101011", 12362 => "0001010100100001", 12363 => "1001001100100001", 12364 => "1110001011111101", 12365 => "1011010100100101", 12366 => "1111111011010001", 12367 => "0100000100110111", 12368 => "0011001110110001", 12369 => "0011010011011100", 12370 => "0101010001100001", 12371 => "1011010001100001", 12372 => "0010111100100111", 12373 => "0000110110010110", 12374 => "1110101110110000", 12375 => "0011010011101001", 12376 => "0010110010010001", 12377 => "0010101101110111", 12378 => "1110101011010111", 12379 => "0000110011011010", 12380 => "1101010111100111", 12381 => "1000111010000101", 12382 => "1110101110101111", 12383 => "0111010011111001", 12384 => "1110111010111110", 12385 => "1011001110000111", 12386 => "1010001011110100", 12387 => "0010000101011011", 12388 => "1101101000011111", 12389 => "0100000110111000", 12390 => "1111111101011100", 12391 => "0010000100000011", 12392 => "1100111111100110", 12393 => "0110010001000110", 12394 => "0111000110101010", 12395 => "1110101010011011", 12396 => "1110001011110100", 12397 => "0001101111110111", 12398 => "1101111001011010", 12399 => "0101111010100010", 12400 => "1000001100010101", 12401 => "1111001000101110", 12402 => "1110010111010111", 12403 => "0111011010100010", 12404 => "1011111010110000", 12405 => "0110010111110100", 12406 => "1101100001001010", 12407 => "1011101010100101", 12408 => "0100100110100110", 12409 => "0010011011001101", 12410 => "0101011001100101", 12411 => "0101011100011000", 12412 => "0110110101101000", 12413 => "0111000010100011", 12414 => "1100000110110001", 12415 => "0011001001100000", 12416 => "0011011111010110", 12417 => "1100100000110111", 12418 => "1100111010000011", 12419 => "0110101010011111", 12420 => "1011011110110101", 12421 => "0111110111011110", 12422 => "1000110111111111", 12423 => "1110010101011110", 12424 => "1100110001100000", 12425 => "1110000001011011", 12426 => "0011100100100011", 12427 => "0000011100000110", 12428 => "0111010110000001", 12429 => "1000010010000110", 12430 => "1101001111000000", 12431 => "0000000110001010", 12432 => "0111001100011101", 12433 => "0110001101010001", 12434 => "1110101010111000", 12435 => "0001101100000010", 12436 => "1110000110001101", 12437 => "1011010110001100", 12438 => "0110000111100111", 12439 => "0101101011010000", 12440 => "1101101010100100", 12441 => "0010111000100111", 12442 => "0101001101100111", 12443 => "1000001101100010", 12444 => "0101111000011010", 12445 => "1110011100011100", 12446 => "1101111101100101", 12447 => "1000111100111100", 12448 => "1001101001011101", 12449 => "1101100001000101", 12450 => "0111011101110110", 12451 => "0100010101000111", 12452 => "1000001100000010", 12453 => "0110000000000101", 12454 => "0001101001101010", 12455 => "1111111110010110", 12456 => "0111101110110101", 12457 => "0010111111010001", 12458 => "1011001101010110", 12459 => "0010011011111010", 12460 => "1100111001110011", 12461 => "0000000000111010", 12462 => "0011110000111000", 12463 => "1110110010011100", 12464 => "0101001100010101", 12465 => "0010101110011000", 12466 => "0100110111000000", 12467 => "1000110010010000", 12468 => "1100100000111000", 12469 => "1011011011000001", 12470 => "1011001000100100", 12471 => "1011011101000101", 12472 => "0101101001000100", 12473 => "1110001110001001", 12474 => "0010010101001011", 12475 => "1011010110100001", 12476 => "1001011011010111", 12477 => "1011010101011101", 12478 => "0011001100110011", 12479 => "1100001011000111", 12480 => "0101111110010100", 12481 => "1100011011100000", 12482 => "0001110101000111", 12483 => "0100111011000111", 12484 => "1101100101011111", 12485 => "1111011000010010", 12486 => "0000110100011011", 12487 => "1100110110000001", 12488 => "1001001101101010", 12489 => "0100010011100111", 12490 => "1011110111000111", 12491 => "0000011100101001", 12492 => "0000011000000001", 12493 => "0111011101100110", 12494 => "0110000110010010", 12495 => "0010000000101010", 12496 => "0011000000110001", 12497 => "0011011000001001", 12498 => "1101101111111110", 12499 => "0010001111001000", 12500 => "1100101100001100", 12501 => "0111001110011000", 12502 => "1100101100111001", 12503 => "1010101100001000", 12504 => "0011111110101001", 12505 => "1100000100101001", 12506 => "1001000101101110", 12507 => "1011101000111101", 12508 => "0100010101011110", 12509 => "1101101001001011", 12510 => "0011111101100010", 12511 => "0101001110110111", 12512 => "0101001010000000", 12513 => "0001011100101001", 12514 => "1100000010000010", 12515 => "1110101110111011", 12516 => "0000011011010100", 12517 => "1101110110110011", 12518 => "0001111010111110", 12519 => "0100110000001110", 12520 => "0000101001011100", 12521 => "1111110100011000", 12522 => "0100011011100110", 12523 => "0010000101100101", 12524 => "0100100000100110", 12525 => "1110011011100010", 12526 => "0001001110000010", 12527 => "1111101110000001", 12528 => "1110010001001001", 12529 => "0101000001011010", 12530 => "0101000111100100", 12531 => "1000010010101011", 12532 => "0100001011111100", 12533 => "1101011011010001", 12534 => "0000001011001100", 12535 => "0111111000111011", 12536 => "1110111110111111", 12537 => "1111100011110101", 12538 => "1011101001001100", 12539 => "1000001110001100", 12540 => "0001000010110110", 12541 => "1010111011010111", 12542 => "0011010101011000", 12543 => "1001010100001000", 12544 => "1011100010110111", 12545 => "0111110001101111", 12546 => "0001000000100111", 12547 => "1101100001011100", 12548 => "1100000000111100", 12549 => "0010111110110101", 12550 => "0000010110000010", 12551 => "1101101011000011", 12552 => "0001000011011111", 12553 => "1001000111110010", 12554 => "1001110010110111", 12555 => "0111001011010010", 12556 => "1000101000011100", 12557 => "0001111110010000", 12558 => "1101100001111011", 12559 => "0001110000001101", 12560 => "1011011011100011", 12561 => "1101011101010000", 12562 => "1111010110100010", 12563 => "0101011000101000", 12564 => "0001110100111011", 12565 => "1100000110000100", 12566 => "1000100000000100", 12567 => "0010001000110001", 12568 => "1111011111001110", 12569 => "1011101111001010", 12570 => "1011001010011011", 12571 => "0100100110000101", 12572 => "0111001110011110", 12573 => "0011000101111111", 12574 => "1101001001010100", 12575 => "1001010100101111", 12576 => "0110011001010101", 12577 => "0100011110101011", 12578 => "1001110010100000", 12579 => "1111010111010001", 12580 => "1010000110001100", 12581 => "0111010000110011", 12582 => "0010110111110101", 12583 => "1010010110010101", 12584 => "1010001110010011", 12585 => "1101110010111010", 12586 => "1110010101000000", 12587 => "1110001001110011", 12588 => "1011100000011000", 12589 => "1100101111010000", 12590 => "0000100101111111", 12591 => "1111101100011000", 12592 => "1000010011000111", 12593 => "1110100111111110", 12594 => "0001111110111010", 12595 => "0100100101100011", 12596 => "1010100000001010", 12597 => "1001110000110011", 12598 => "1010101001111000", 12599 => "0001010100100011", 12600 => "0110110101011110", 12601 => "1010001000010001", 12602 => "0110000111101010", 12603 => "1100101000101101", 12604 => "0101110011000011", 12605 => "1111110111101110", 12606 => "1100110101101000", 12607 => "0110000111010010", 12608 => "1000011010010011", 12609 => "1100100001111010", 12610 => "1100101000101110", 12611 => "1011010010000101", 12612 => "1000011010110100", 12613 => "1101100111010001", 12614 => "0111111010001010", 12615 => "0000110011111100", 12616 => "1111000001101101", 12617 => "0100110101100101", 12618 => "1000101001100011", 12619 => "1101110010001100", 12620 => "1001000101100010", 12621 => "1001000011011101", 12622 => "0011111111110100", 12623 => "0010111101010111", 12624 => "1100010011100101", 12625 => "1001011011001111", 12626 => "1100111010100010", 12627 => "0000100100010110", 12628 => "0010010000010101", 12629 => "0000110101101101", 12630 => "1001111011001110", 12631 => "1110011010100000", 12632 => "0000011000100100", 12633 => "0000000110100000", 12634 => "0110101001010100", 12635 => "1110001001010000", 12636 => "0000001000001100", 12637 => "0010110011100011", 12638 => "1100100000011001", 12639 => "0100001001111110", 12640 => "1010000010101111", 12641 => "1101011111010100", 12642 => "0110110110111111", 12643 => "1101010011101100", 12644 => "0101110100110110", 12645 => "0000001100001011", 12646 => "1101111011100110", 12647 => "0010110100011100", 12648 => "1001000110101001", 12649 => "1110111110011101", 12650 => "1111101010001100", 12651 => "1101011100110110", 12652 => "0100110011010100", 12653 => "0100101101110011", 12654 => "1101111111111110", 12655 => "0011000000001100", 12656 => "1000001011110010", 12657 => "1010011101101000", 12658 => "1001100100011011", 12659 => "1011110101011101", 12660 => "1111101100000111", 12661 => "1100000001110011", 12662 => "0101110100000010", 12663 => "1000100010111110", 12664 => "1101111000010110", 12665 => "1001110100010101", 12666 => "1000110000100110", 12667 => "1001100110111101", 12668 => "0011100100010111", 12669 => "0001001110101100", 12670 => "0101101110000100", 12671 => "0100000101110101", 12672 => "0101011100011100", 12673 => "1100111100000110", 12674 => "1010001101001100", 12675 => "0101010000100001", 12676 => "1111011101001111", 12677 => "1111101100111100", 12678 => "1000110101101011", 12679 => "0001110110100011", 12680 => "1110001000000101", 12681 => "0110111001101100", 12682 => "0110010100000101", 12683 => "0110001101111000", 12684 => "1010110110100000", 12685 => "1011001110001011", 12686 => "1000100110001100", 12687 => "0100001101101000", 12688 => "0011000111000101", 12689 => "1000101010001001", 12690 => "1000101110101111", 12691 => "0100001001100000", 12692 => "1001010000010001", 12693 => "0110100001010110", 12694 => "1100000001010111", 12695 => "1111010011100001", 12696 => "1100011011011010", 12697 => "0110000101001001", 12698 => "1111111110000101", 12699 => "0010100111000100", 12700 => "1110000011010100", 12701 => "0010110110010010", 12702 => "0001011000100111", 12703 => "0110001011000100", 12704 => "1101110110001101", 12705 => "1000010100101100", 12706 => "0010110001110110", 12707 => "1010001110110100", 12708 => "0101010111001010", 12709 => "1110111011110110", 12710 => "0110000000101010", 12711 => "0011010000001110", 12712 => "0111111101111000", 12713 => "1100100111100100", 12714 => "1011111101000111", 12715 => "0101000100111100", 12716 => "1100111110111101", 12717 => "0110100011010001", 12718 => "0000011010000101", 12719 => "0011110011011001", 12720 => "1111001101001100", 12721 => "0001111100001101", 12722 => "0111010000011010", 12723 => "1001101111101001", 12724 => "0111011010111011", 12725 => "0000100010101100", 12726 => "0010101011111100", 12727 => "1001100010100000", 12728 => "0110010100011111", 12729 => "1011010010000101", 12730 => "1011000101100000", 12731 => "0001111011011111", 12732 => "1110101000100001", 12733 => "1100010011110101", 12734 => "0010010001101010", 12735 => "1010011010010010", 12736 => "1000001010011100", 12737 => "1011001000011001", 12738 => "0111010010110111", 12739 => "1101011100011010", 12740 => "1101110110010111", 12741 => "1000000100001111", 12742 => "1000101010101101", 12743 => "1001011111110000", 12744 => "1110110111000110", 12745 => "1110100110001110", 12746 => "1001001011011011", 12747 => "0011111011010011", 12748 => "1001000111001110", 12749 => "0001100110011011", 12750 => "0101110010100100", 12751 => "1110001010000110", 12752 => "1110100100001001", 12753 => "0011100110110111", 12754 => "0111001010001100", 12755 => "1010110101110000", 12756 => "0000100001101100", 12757 => "1001000110001010", 12758 => "0010101110000001", 12759 => "0001110010011111", 12760 => "0100100010100101", 12761 => "0011110101110101", 12762 => "1110110101110110", 12763 => "1111100111001011", 12764 => "1111010111101010", 12765 => "0111110010010111", 12766 => "0000010001100001", 12767 => "0110100011100000", 12768 => "1110111001011100", 12769 => "1110110001101011", 12770 => "1110000101110000", 12771 => "0011100001100111", 12772 => "1101010010101100", 12773 => "1000001001000101", 12774 => "0111101001101101", 12775 => "1000111010000011", 12776 => "1010111010001010", 12777 => "1010111101101111", 12778 => "0010010110100010", 12779 => "0010100110100000", 12780 => "1000001010011000", 12781 => "0000011101011110", 12782 => "1111000010111001", 12783 => "1010011001010011", 12784 => "1001001011101100", 12785 => "0100001000001001", 12786 => "1001111000110001", 12787 => "1110011000111010", 12788 => "0110000111100110", 12789 => "0100101100000001", 12790 => "0101000001110011", 12791 => "1000110000110011", 12792 => "0010001001101011", 12793 => "0111011001010000", 12794 => "0011011110111000", 12795 => "1100110101000101", 12796 => "1000011100010111", 12797 => "0000101010000010", 12798 => "1100111000100011", 12799 => "0100100110111011", 12800 => "1101110001101111", 12801 => "1110010100000111", 12802 => "0100011011000110", 12803 => "0010110000111000", 12804 => "0000000001010111", 12805 => "0000000101010110", 12806 => "1000011010100010", 12807 => "1111100010101110", 12808 => "0001111010010111", 12809 => "1001000110001000", 12810 => "0111011111010010", 12811 => "0001110001111101", 12812 => "1101101001111101", 12813 => "1011011111010010", 12814 => "0111111100111000", 12815 => "0000010011111001", 12816 => "1000101110000100", 12817 => "0000010010100101", 12818 => "0110101100100101", 12819 => "1110011000011011", 12820 => "0001100110001111", 12821 => "0011010010001001", 12822 => "0100110110000001", 12823 => "0000101001110111", 12824 => "1010100011011110", 12825 => "0001101100101000", 12826 => "1101001001000000", 12827 => "1111011011010101", 12828 => "0111111100011010", 12829 => "1110001101100111", 12830 => "1100110010111111", 12831 => "1100100111000101", 12832 => "0101010100000010", 12833 => "0001111111101111", 12834 => "1000000100001011", 12835 => "1100000101111011", 12836 => "0010001111111101", 12837 => "1000110111001100", 12838 => "1000101011101100", 12839 => "1010111000010001", 12840 => "0101011111111101", 12841 => "0010011111100111", 12842 => "0111010000011000", 12843 => "1001110000010110", 12844 => "1110001100110000", 12845 => "1110101000010011", 12846 => "1011001001110111", 12847 => "1000111101100101", 12848 => "1011001011100100", 12849 => "1011010001000000", 12850 => "0110011100111101", 12851 => "1111010100010100", 12852 => "0000110100011010", 12853 => "0000111110010110", 12854 => "0010000001100000", 12855 => "1001010100110010", 12856 => "1110101010110011", 12857 => "0000011011010000", 12858 => "0011100001111010", 12859 => "0101100000111011", 12860 => "0101110011101011", 12861 => "0110101000010111", 12862 => "1000011000000011", 12863 => "0010100110101001", 12864 => "1111010100100101", 12865 => "0100001001011111", 12866 => "1110101100101110", 12867 => "1011111100110010", 12868 => "0011100100000101", 12869 => "0011001110001100", 12870 => "1000100010010101", 12871 => "1101011010010101", 12872 => "1000101000010100", 12873 => "1111101011101010", 12874 => "0110010111001011", 12875 => "1010011010001101", 12876 => "0101011000000110", 12877 => "1111111011111011", 12878 => "0000001100001100", 12879 => "1000100101011110", 12880 => "1001000010101110", 12881 => "0100001001010001", 12882 => "0011111110111010", 12883 => "0010010010110111", 12884 => "1000100000100110", 12885 => "1100011110001101", 12886 => "1001001111010010", 12887 => "0100011111110111", 12888 => "1011101101110100", 12889 => "0011010110100100", 12890 => "0101101101101010", 12891 => "0101010001101100", 12892 => "1010100100100000", 12893 => "0100110010110111", 12894 => "0110101101011010", 12895 => "1001000110001110", 12896 => "1101101001001101", 12897 => "0001100001100100", 12898 => "0011001110101000", 12899 => "0100100111101100", 12900 => "0100011101000000", 12901 => "0011101011110101", 12902 => "0011000000110001", 12903 => "0011111100101101", 12904 => "0111000011100111", 12905 => "0111111001010011", 12906 => "0001110110011010", 12907 => "1010000001100011", 12908 => "1010000000001101", 12909 => "0000011010110001", 12910 => "1000111101000000", 12911 => "1101001011111100", 12912 => "0010100110000011", 12913 => "1110101101101001", 12914 => "1100000110011101", 12915 => "0001001000110100", 12916 => "1010111010011000", 12917 => "1001000000100000", 12918 => "0011010000101001", 12919 => "0011101000001100", 12920 => "1101111010001000", 12921 => "0001000101110101", 12922 => "1000110101100101", 12923 => "0111001111101011", 12924 => "0111101101010011", 12925 => "0001010111010110", 12926 => "1011111000010101", 12927 => "0011000000110110", 12928 => "1100111011101101", 12929 => "0101100011011110", 12930 => "1001100001000111", 12931 => "1110001101001110", 12932 => "1100100110111011", 12933 => "0000000110011010", 12934 => "1001111011011100", 12935 => "1000011010001100", 12936 => "0001001111110010", 12937 => "0100101001110111", 12938 => "1010101111011001", 12939 => "1111101001010110", 12940 => "0011011010011001", 12941 => "0000100000001100", 12942 => "0111011110100110", 12943 => "0110100011111000", 12944 => "1100110100110110", 12945 => "0111101001110111", 12946 => "1001001010010111", 12947 => "1010011100011111", 12948 => "0010000001111101", 12949 => "1010010100100010", 12950 => "0111101111010011", 12951 => "0100111111001110", 12952 => "0000100110100011", 12953 => "0100101110011111", 12954 => "0111001110001110", 12955 => "1110000010100010", 12956 => "1000101011000011", 12957 => "1001111110011000", 12958 => "0100011100000000", 12959 => "0000100000101110", 12960 => "0000101001010111", 12961 => "0100100010011101", 12962 => "1000100010110010", 12963 => "0000110111101100", 12964 => "1010001100111110", 12965 => "1000100100101111", 12966 => "0000100101001100", 12967 => "1011011111011100", 12968 => "1011101101101111", 12969 => "1011010011000100", 12970 => "0010000110001011", 12971 => "0101001110110110", 12972 => "0000110110110101", 12973 => "1110001001100101", 12974 => "0010010011100000", 12975 => "1101011000100110", 12976 => "1001000111110100", 12977 => "1101100010111111", 12978 => "1000001101111001", 12979 => "1111110101100100", 12980 => "1011011010001001", 12981 => "0001000011011110", 12982 => "0100010110100100", 12983 => "0101010011001010", 12984 => "0100111110100000", 12985 => "0010101101100000", 12986 => "0101111110100101", 12987 => "0101100111110010", 12988 => "1010001111011011", 12989 => "1011000010000100", 12990 => "0011000110011110", 12991 => "0101100000111010", 12992 => "1000111111101100", 12993 => "0000011100110111", 12994 => "1110110111110111", 12995 => "0010011010000111", 12996 => "1010111010110100", 12997 => "0100111000111001", 12998 => "1111011000111110", 12999 => "1001101010000101", 13000 => "1110011110101101", 13001 => "1111011010110010", 13002 => "1001111001101000", 13003 => "0101011001101010", 13004 => "1011111001100001", 13005 => "0110000100001110", 13006 => "1001001010111001", 13007 => "0000110011011000", 13008 => "1100010000110000", 13009 => "0100010000100010", 13010 => "0010100010101010", 13011 => "1111110010111001", 13012 => "1101010010011010", 13013 => "1100011110011010", 13014 => "1001111010001010", 13015 => "1010111000000101", 13016 => "1101010001011111", 13017 => "0000100110011000", 13018 => "0101011100100100", 13019 => "1011110111000110", 13020 => "1100011001010110", 13021 => "0010110111111110", 13022 => "0000001011011111", 13023 => "0001000101110111", 13024 => "0011111111000111", 13025 => "0001011000010111", 13026 => "1101100010000001", 13027 => "0000110110001010", 13028 => "1001010101110100", 13029 => "1011001001010100", 13030 => "0101111001110101", 13031 => "1011000010111000", 13032 => "0100101010110000", 13033 => "0001101111001111", 13034 => "1111011111001101", 13035 => "1100001001000001", 13036 => "0101101000110110", 13037 => "1011010010000110", 13038 => "0011101001000110", 13039 => "0001001100110001", 13040 => "1000100101110100", 13041 => "1000011000101100", 13042 => "1110100010100000", 13043 => "0010110101000100", 13044 => "1110010110001101", 13045 => "0101110100110010", 13046 => "0000101110101010", 13047 => "1000111100011000", 13048 => "1011000100110001", 13049 => "0000011000110000", 13050 => "1010111111011011", 13051 => "0111011101110011", 13052 => "1100100101010110", 13053 => "1101001111101010", 13054 => "1001000001001001", 13055 => "1101111111110111", 13056 => "0011101011101010", 13057 => "0111100101000010", 13058 => "0111001100000000", 13059 => "1001011110001001", 13060 => "0111001101111010", 13061 => "0100110000010110", 13062 => "0010000110101010", 13063 => "1100101010011001", 13064 => "0000001010001011", 13065 => "1001011110110000", 13066 => "0011001000000000", 13067 => "1100011101110011", 13068 => "1101000011011001", 13069 => "0001100001110101", 13070 => "1010111101011111", 13071 => "1111010110101100", 13072 => "0000111111110111", 13073 => "0011101100010110", 13074 => "1010101010111000", 13075 => "0101100110101110", 13076 => "0100011101101001", 13077 => "1111010010000010", 13078 => "1001010101010110", 13079 => "1010001100010011", 13080 => "1100100101000110", 13081 => "1111101001000110", 13082 => "1000101110010011", 13083 => "0100011001011000", 13084 => "1010110110111000", 13085 => "0010001101111100", 13086 => "1100011110110100", 13087 => "1110011110110110", 13088 => "0111001010010100", 13089 => "0011001000000110", 13090 => "1110011010111100", 13091 => "1101101011011001", 13092 => "1101000000011101", 13093 => "1000110100011101", 13094 => "1001000100011011", 13095 => "1000000001111100", 13096 => "0011010110011110", 13097 => "0011001001001101", 13098 => "0011001100101000", 13099 => "1000100101010101", 13100 => "0110011111010011", 13101 => "0011011111011001", 13102 => "0010110110101001", 13103 => "1110101011101111", 13104 => "1101001001110011", 13105 => "0010100000111000", 13106 => "1110101111111001", 13107 => "1101110000101001", 13108 => "0000111101100101", 13109 => "0100010001111101", 13110 => "1101010111010110", 13111 => "1000111001101111", 13112 => "0001111010000000", 13113 => "1111100001000011", 13114 => "0111000110011010", 13115 => "0110110111100011", 13116 => "0101000001011010", 13117 => "1000110101011011", 13118 => "1000110010110110", 13119 => "1011010000011101", 13120 => "1110110100110001", 13121 => "1011101100101110", 13122 => "1001001001000110", 13123 => "0111111010001101", 13124 => "1000001101110000", 13125 => "1100011110000111", 13126 => "0100100101111010", 13127 => "0010101011101011", 13128 => "1110011100000010", 13129 => "0000000100101001", 13130 => "1101100111010001", 13131 => "0000110000010010", 13132 => "0000100010111011", 13133 => "1000100000111010", 13134 => "0011110100010011", 13135 => "1011011001011101", 13136 => "1010100111001011", 13137 => "0111101010000100", 13138 => "1100111000001111", 13139 => "1000101111100101", 13140 => "1110111010100011", 13141 => "0001000110110111", 13142 => "0001011111110111", 13143 => "0101000010001010", 13144 => "0000011011111100", 13145 => "1011001111010110", 13146 => "0001001010011101", 13147 => "0101100101110001", 13148 => "1000010010100110", 13149 => "0100111011100111", 13150 => "1000101010100001", 13151 => "1000101111101101", 13152 => "1001100010001011", 13153 => "1111101010010011", 13154 => "0110100001010011", 13155 => "0010010011110011", 13156 => "0001101000110111", 13157 => "1010110100100010", 13158 => "1010110000010111", 13159 => "1001101110000001", 13160 => "0001001010110110", 13161 => "0111011001111111", 13162 => "0011100110001001", 13163 => "0010110001000110", 13164 => "1001101111001100", 13165 => "0011010011110100", 13166 => "1110100010001100", 13167 => "1101111001110001", 13168 => "0110000001000011", 13169 => "1111100101010111", 13170 => "1110111001100110", 13171 => "0000100110011111", 13172 => "1011010111110000", 13173 => "1101011110111010", 13174 => "1000101011111110", 13175 => "1101110110010001", 13176 => "1011010110100101", 13177 => "0010111110100001", 13178 => "1100011110111111", 13179 => "1110001010110100", 13180 => "0100110001111111", 13181 => "1111010110101010", 13182 => "0001010001111100", 13183 => "0001000011001100", 13184 => "0101110111000001", 13185 => "0000101101111110", 13186 => "1100101001000001", 13187 => "0100110111010100", 13188 => "1011110100110000", 13189 => "0101011100100010", 13190 => "1010111111110010", 13191 => "1000010001001011", 13192 => "1000110100100111", 13193 => "0100011100101100", 13194 => "1111110011001110", 13195 => "0010011100011010", 13196 => "0010000001001100", 13197 => "0010011100110101", 13198 => "1000001000101110", 13199 => "0000000001010100", 13200 => "0101010110011000", 13201 => "1101000110010101", 13202 => "0110101010101100", 13203 => "1010001000000110", 13204 => "0111110110111000", 13205 => "0010110100010101", 13206 => "1001010100000110", 13207 => "0101101101011010", 13208 => "0011011000100011", 13209 => "1110000111000101", 13210 => "1010011101101110", 13211 => "0110011100010000", 13212 => "1010001000000111", 13213 => "1011111100011001", 13214 => "0010001101100001", 13215 => "1111100100010000", 13216 => "1101110000100010", 13217 => "0100100110001000", 13218 => "1101111000101001", 13219 => "0010111001010111", 13220 => "0101101111011011", 13221 => "0110101111111110", 13222 => "0010000110100010", 13223 => "0111110110011000", 13224 => "0001111110010011", 13225 => "0111111001110100", 13226 => "1111100101011000", 13227 => "0111111000101110", 13228 => "1001011100000110", 13229 => "0100001101101110", 13230 => "0001001010010000", 13231 => "1111000001000001", 13232 => "0100001001100011", 13233 => "0011101110111011", 13234 => "0110110100110101", 13235 => "0001100011111010", 13236 => "1111000000010100", 13237 => "0110110000111110", 13238 => "1011011111001010", 13239 => "0110111001101110", 13240 => "0110010000110110", 13241 => "1111111000110101", 13242 => "1011110110011100", 13243 => "0001101111001101", 13244 => "0001010001011111", 13245 => "0101110100011001", 13246 => "0101100100011100", 13247 => "0101110111000010", 13248 => "1110111111110100", 13249 => "0111100100111110", 13250 => "1110111101000011", 13251 => "0101100100110010", 13252 => "0001100010010000", 13253 => "1101101100001010", 13254 => "0001010011010010", 13255 => "0000010000001001", 13256 => "0100111110110100", 13257 => "0000110111101011", 13258 => "1100011010010110", 13259 => "0110101110000101", 13260 => "0011110001110010", 13261 => "0100000011101000", 13262 => "1000111100000000", 13263 => "0111011011001110", 13264 => "1111011111001100", 13265 => "1010010111011010", 13266 => "0110100000101000", 13267 => "1111000101101111", 13268 => "0111000011011110", 13269 => "0001011101010110", 13270 => "1111001110100000", 13271 => "0010011101001000", 13272 => "0011110100011011", 13273 => "0110101011000111", 13274 => "0000000011101011", 13275 => "1011000001010010", 13276 => "0111100101100100", 13277 => "1101100111010000", 13278 => "1001110111011111", 13279 => "1010111110100100", 13280 => "1001000001111101", 13281 => "0111000110010101", 13282 => "1110011010101011", 13283 => "1100001010001011", 13284 => "0001001011100101", 13285 => "0001001011100100", 13286 => "1111101111010001", 13287 => "1011001010110100", 13288 => "0110010111010011", 13289 => "0010001100100111", 13290 => "0111110000111110", 13291 => "1000101011111100", 13292 => "0110010100110001", 13293 => "0011110100111100", 13294 => "0111100100110010", 13295 => "1110101001001100", 13296 => "0001010110000000", 13297 => "0000111111011001", 13298 => "0111100001100110", 13299 => "0010000110000010", 13300 => "0101010010110001", 13301 => "0100010000110011", 13302 => "0100000010111011", 13303 => "0110101000110110", 13304 => "1110000100001011", 13305 => "0100110001100001", 13306 => "1110001001111001", 13307 => "0100010111011111", 13308 => "1110100101011101", 13309 => "0001001011001000", 13310 => "0100000110101110", 13311 => "0110100001110110", 13312 => "1010010001010101", 13313 => "1101011000111010", 13314 => "0000110101011110", 13315 => "0101110101010000", 13316 => "1101110011001010", 13317 => "0110100000100101", 13318 => "0111010011100110", 13319 => "0011010110100101", 13320 => "1011110011101011", 13321 => "0011101100001000", 13322 => "0000100111001000", 13323 => "0000000101010101", 13324 => "0111011001111110", 13325 => "1110111101101110", 13326 => "1000000110001010", 13327 => "1001001011100100", 13328 => "0011111000111111", 13329 => "0001101110101101", 13330 => "1101011111101011", 13331 => "0100101101011010", 13332 => "0000111001011000", 13333 => "1011010010111011", 13334 => "0101100000111100", 13335 => "1100010011101000", 13336 => "0011010011011110", 13337 => "0000111100000010", 13338 => "1011000010110110", 13339 => "1001110101100010", 13340 => "1001000010111011", 13341 => "0010001011110011", 13342 => "0101011110001111", 13343 => "1011010110011001", 13344 => "0110010111000101", 13345 => "1110110101100110", 13346 => "0100000110111000", 13347 => "0110011101000000", 13348 => "1000000110000001", 13349 => "1111001001110011", 13350 => "1011000011100100", 13351 => "1011010010110111", 13352 => "0101111100110011", 13353 => "1011110010110001", 13354 => "1000110000011101", 13355 => "0111010010110010", 13356 => "1100110101110110", 13357 => "1110001101100111", 13358 => "1000001000011011", 13359 => "1010000100110010", 13360 => "0001110110111101", 13361 => "0101011100010011", 13362 => "0110111100110011", 13363 => "1110100001101101", 13364 => "0100001101010100", 13365 => "0100101111100001", 13366 => "0100110100001100", 13367 => "0001001010111100", 13368 => "0011000101010101", 13369 => "0000001101101010", 13370 => "1101110110001011", 13371 => "0100100011010010", 13372 => "1011110000011010", 13373 => "0110101110011101", 13374 => "1010000011010100", 13375 => "0011110011001011", 13376 => "0011111000110011", 13377 => "0100110101101101", 13378 => "0101111101001101", 13379 => "1001111011101100", 13380 => "0110010000100011", 13381 => "0010110001100011", 13382 => "0101100111110100", 13383 => "1010011011001010", 13384 => "1001011011100101", 13385 => "1011111011101000", 13386 => "1110000101111101", 13387 => "1001100111101010", 13388 => "0000111110000011", 13389 => "1100011110011000", 13390 => "1111111100110000", 13391 => "1010111100010111", 13392 => "1010000001100010", 13393 => "0000111000111111", 13394 => "0000110000011110", 13395 => "0100000011001101", 13396 => "0110101101101001", 13397 => "1011011110100001", 13398 => "1100000101010100", 13399 => "0100110100111000", 13400 => "0100000010010001", 13401 => "1011000011110001", 13402 => "0000010101111110", 13403 => "1000000001101010", 13404 => "0100111001011111", 13405 => "0001000100001110", 13406 => "1100010110011110", 13407 => "0101001110010101", 13408 => "0100011001110101", 13409 => "0100010111010100", 13410 => "0111000010011001", 13411 => "1111011110001001", 13412 => "1110011100100000", 13413 => "1100101110001010", 13414 => "1110100100101010", 13415 => "1001100110101100", 13416 => "0111110101110111", 13417 => "1001000111111101", 13418 => "1011000001111011", 13419 => "1001000010011100", 13420 => "0000111111011100", 13421 => "0110001111101101", 13422 => "1000111001000010", 13423 => "0101011111110101", 13424 => "0110111001010010", 13425 => "1101001100100001", 13426 => "0110101101000110", 13427 => "0001001010101001", 13428 => "0001010001011110", 13429 => "1000011100000111", 13430 => "1000101000010100", 13431 => "1101111010110111", 13432 => "0101111100100011", 13433 => "1110010110111000", 13434 => "1011111101101110", 13435 => "0010101110100100", 13436 => "1010100010101010", 13437 => "1001101101101101", 13438 => "1001110000001100", 13439 => "0010011101010110", 13440 => "0110010111101101", 13441 => "0001000010100110", 13442 => "1010110100000101", 13443 => "0011011011100110", 13444 => "1101100011100011", 13445 => "1111111110110111", 13446 => "0100011100110000", 13447 => "0101111011011000", 13448 => "0000111010000101", 13449 => "0001110011011001", 13450 => "0010010011110000", 13451 => "1110101101011010", 13452 => "1000011001000001", 13453 => "1110011010011011", 13454 => "1110100000001010", 13455 => "0001011111010110", 13456 => "1110101000011000", 13457 => "1110011111010100", 13458 => "1100101111110110", 13459 => "0011010000010011", 13460 => "0000101011111011", 13461 => "0000010101000111", 13462 => "0111110100001001", 13463 => "0110110001011110", 13464 => "0010110000101110", 13465 => "1001110111000110", 13466 => "1101100001110010", 13467 => "0101111001110111", 13468 => "1110011111011001", 13469 => "0000010010110110", 13470 => "0110001100101101", 13471 => "0100001000000001", 13472 => "1000000111110010", 13473 => "1110001011101111", 13474 => "0000110110111111", 13475 => "1001001001011110", 13476 => "0001000010010100", 13477 => "1000110011011110", 13478 => "0110010110000001", 13479 => "0001011110011111", 13480 => "1001001010010100", 13481 => "1100111101000011", 13482 => "0101001010111011", 13483 => "0001000101001000", 13484 => "0010110111001000", 13485 => "1110010000011001", 13486 => "0011010111000010", 13487 => "1001110100100001", 13488 => "1011101101100100", 13489 => "1001011101110011", 13490 => "0001000100011011", 13491 => "0101100010011001", 13492 => "1111001100010101", 13493 => "1001100111001110", 13494 => "0000000100000101", 13495 => "1001010000010101", 13496 => "1010101110111100", 13497 => "0011001111001011", 13498 => "1010110101111110", 13499 => "0101111111101111", 13500 => "1100100010000101", 13501 => "0111101001101100", 13502 => "1110000100101000", 13503 => "0000111010000010", 13504 => "0011110001100100", 13505 => "0011011010101111", 13506 => "0001100111000101", 13507 => "0100110001100100", 13508 => "1001001011110101", 13509 => "0110010110101011", 13510 => "1101000101100111", 13511 => "1110100111000000", 13512 => "1011000101100011", 13513 => "0001111101001111", 13514 => "1000000011111001", 13515 => "0010010101011001", 13516 => "0001111011001111", 13517 => "1001110000110010", 13518 => "1111011010010100", 13519 => "1001110001110011", 13520 => "1100111111001000", 13521 => "0110000111111100", 13522 => "1110110011110011", 13523 => "1010111101100101", 13524 => "1110110010100000", 13525 => "0000110100011100", 13526 => "1011100000001000", 13527 => "1010101101111000", 13528 => "1000111010101111", 13529 => "0010100100011000", 13530 => "1011101111011111", 13531 => "0100001011110100", 13532 => "1010110111100101", 13533 => "0010010111011101", 13534 => "0011011100100011", 13535 => "0000111100111101", 13536 => "0001111001011000", 13537 => "0110011010101000", 13538 => "1111110001001111", 13539 => "1001010111000111", 13540 => "1100101100100110", 13541 => "0000111001001111", 13542 => "0101100101001001", 13543 => "0101001101111100", 13544 => "0001011111111001", 13545 => "1110011000101001", 13546 => "0111100001011010", 13547 => "1111111010010001", 13548 => "0111101010010101", 13549 => "0001000101110001", 13550 => "1101101001100011", 13551 => "0111111101010011", 13552 => "1001010101011001", 13553 => "1001101011101100", 13554 => "1100111010001011", 13555 => "1010100000110010", 13556 => "0001101000010111", 13557 => "1100110101010000", 13558 => "0010100101001100", 13559 => "0011011110010100", 13560 => "1000010111001001", 13561 => "1101000000011001", 13562 => "1111011010011001", 13563 => "0100100011010010", 13564 => "1100001001100101", 13565 => "0100001001110011", 13566 => "1110110001101001", 13567 => "1111110000010100", 13568 => "0111110001101110", 13569 => "1101000110011100", 13570 => "0110001011111100", 13571 => "1010001101101101", 13572 => "0011010000011101", 13573 => "1100111011101110", 13574 => "1000011000011100", 13575 => "0110101000100100", 13576 => "1110011100100000", 13577 => "1011101101101001", 13578 => "1110010011110000", 13579 => "0100001010010110", 13580 => "0010110010011111", 13581 => "0100011101011111", 13582 => "0000011100110010", 13583 => "1111011110110010", 13584 => "0000110101000110", 13585 => "0110110010011101", 13586 => "1010110001010001", 13587 => "1100110000100100", 13588 => "1101001110101001", 13589 => "0110100110100111", 13590 => "0000101000101010", 13591 => "1001011111101110", 13592 => "1110110101000011", 13593 => "1110010001111110", 13594 => "0000011001010110", 13595 => "1000101101111001", 13596 => "1110100011110111", 13597 => "1110111000001011", 13598 => "0000110010000010", 13599 => "0011011100010001", 13600 => "1011000101011101", 13601 => "0011111111011111", 13602 => "0001110001000101", 13603 => "1101011000111100", 13604 => "1010110011001010", 13605 => "0011001000010110", 13606 => "1100001110011001", 13607 => "0110000110101101", 13608 => "0001000001111001", 13609 => "1111111010010100", 13610 => "1011101111001110", 13611 => "0001010000100000", 13612 => "1010110011001001", 13613 => "1010101010100001", 13614 => "1000000111110000", 13615 => "0011010010011001", 13616 => "1101111001011111", 13617 => "1010001011110011", 13618 => "1111101001001001", 13619 => "1000010100111001", 13620 => "1000111001110001", 13621 => "0001101000101010", 13622 => "0111000100101001", 13623 => "0000101101111111", 13624 => "0001011011011000", 13625 => "0010110000011010", 13626 => "0110011100110011", 13627 => "1010010100100010", 13628 => "0001010011011011", 13629 => "1101010100010001", 13630 => "1110111011101101", 13631 => "0100011111010110", 13632 => "1100101011110110", 13633 => "0001100001111101", 13634 => "0110011011000000", 13635 => "0010010101100011", 13636 => "1011010110110000", 13637 => "0011111110110000", 13638 => "1010101110111111", 13639 => "0111011101111010", 13640 => "1011110100111010", 13641 => "0001011110101100", 13642 => "1000100000001000", 13643 => "1111011100011111", 13644 => "1110101000100010", 13645 => "0010100000001100", 13646 => "0111101000010011", 13647 => "1001100010001010", 13648 => "1110011001110010", 13649 => "1010011010010111", 13650 => "0110011010011101", 13651 => "1111110111101111", 13652 => "0000101101110111", 13653 => "1110010011000001", 13654 => "1010101110111001", 13655 => "0011100100111101", 13656 => "1001010110111011", 13657 => "0110101011100101", 13658 => "1001110101010110", 13659 => "1000010110011010", 13660 => "1000001010001000", 13661 => "0001100101001011", 13662 => "0011100111001000", 13663 => "1110110001000011", 13664 => "0111111001010000", 13665 => "1001000111100110", 13666 => "1111001100110101", 13667 => "0011000001000101", 13668 => "1100100100110011", 13669 => "0001100110000100", 13670 => "1011011101000011", 13671 => "0100110001011101", 13672 => "0010101100111100", 13673 => "1001001111100011", 13674 => "0101111101001010", 13675 => "1111011101110101", 13676 => "0010010101001011", 13677 => "0010010101010001", 13678 => "0010001001111110", 13679 => "0111100000100111", 13680 => "0100000111110101", 13681 => "0111000101100111", 13682 => "1001001110010011", 13683 => "1000011010000110", 13684 => "0111110100001010", 13685 => "0110000000100110", 13686 => "0000111111010011", 13687 => "1001110100110111", 13688 => "1100111010010001", 13689 => "0010011110000101", 13690 => "0100000010000111", 13691 => "0010111000000101", 13692 => "1111101111010110", 13693 => "1001011010110000", 13694 => "1111010001011010", 13695 => "0001011111010000", 13696 => "1001011010010110", 13697 => "0001001001100110", 13698 => "0001110000111110", 13699 => "1101001110101001", 13700 => "0101110000000011", 13701 => "0100100000100000", 13702 => "0100111100111110", 13703 => "0111000010011100", 13704 => "0101001101010010", 13705 => "0111011010010001", 13706 => "1100001000000011", 13707 => "1100011010000110", 13708 => "1100010111101010", 13709 => "0101010010001100", 13710 => "0110100101110100", 13711 => "1001111011111011", 13712 => "0101011110010011", 13713 => "0111001000010001", 13714 => "1100100000110000", 13715 => "0111110110011010", 13716 => "0100111110101000", 13717 => "0001110001000011", 13718 => "0100001101001111", 13719 => "0000100110010100", 13720 => "1110110001010000", 13721 => "1001111011000010", 13722 => "1000010010110001", 13723 => "1101010100001111", 13724 => "0000001111111011", 13725 => "1101110111101100", 13726 => "1011000110001011", 13727 => "1101010110010100", 13728 => "0010100001100111", 13729 => "1110111001010000", 13730 => "1101110110110100", 13731 => "0011111010110000", 13732 => "0001110010001000", 13733 => "0010100101011110", 13734 => "1100111011101100", 13735 => "0100111010011100", 13736 => "1010011100111001", 13737 => "1000001011100111", 13738 => "1011110111011111", 13739 => "0111000011101110", 13740 => "0010110000000000", 13741 => "1101000011111001", 13742 => "1100011000111000", 13743 => "0101011110111011", 13744 => "1101001111000000", 13745 => "1110100101100101", 13746 => "1010111011111101", 13747 => "1010010100001100", 13748 => "0011111110110011", 13749 => "0100100110111011", 13750 => "1000111010111111", 13751 => "0011101011000110", 13752 => "1010111001111100", 13753 => "1001001010101000", 13754 => "1000010001111111", 13755 => "0010111001011111", 13756 => "0000101101000101", 13757 => "1100011001000011", 13758 => "0001000110010110", 13759 => "1011101010001001", 13760 => "1000100101011000", 13761 => "1100101010010000", 13762 => "1111111101001101", 13763 => "1111010111101000", 13764 => "0111011001101010", 13765 => "1010001111010000", 13766 => "1000000010100001", 13767 => "1100110011011001", 13768 => "1011100110100011", 13769 => "0111110110001000", 13770 => "0110110111010111", 13771 => "0111001110110101", 13772 => "1010111010110101", 13773 => "0000101010000101", 13774 => "0010010100010011", 13775 => "1000100100100111", 13776 => "1101111111011111", 13777 => "1010011001000001", 13778 => "1111011000100110", 13779 => "1100001000101111", 13780 => "1001101110111011", 13781 => "0111010100111100", 13782 => "0101111110000110", 13783 => "0001010000101110", 13784 => "1000100001110001", 13785 => "0110000010010010", 13786 => "0110101110111000", 13787 => "1111110111111101", 13788 => "1000011111010010", 13789 => "0010110000000100", 13790 => "1111001000000100", 13791 => "1000001010001101", 13792 => "0001101111100001", 13793 => "0111100011011111", 13794 => "0010000001001101", 13795 => "1000001111111001", 13796 => "1111001000000001", 13797 => "0100000010110001", 13798 => "1111011101101011", 13799 => "1001000111010001", 13800 => "0101111000001010", 13801 => "0110100100010010", 13802 => "1011011101001100", 13803 => "1100011111010101", 13804 => "0110100010100111", 13805 => "1011101000110100", 13806 => "1110000101111110", 13807 => "0111000111111110", 13808 => "1001001010011100", 13809 => "1011110000110111", 13810 => "0000001101011010", 13811 => "0010110111011101", 13812 => "0011111011111011", 13813 => "0011100111001110", 13814 => "1111100111011000", 13815 => "0100011000111100", 13816 => "0000011011001100", 13817 => "1101110111000110", 13818 => "0111111011010010", 13819 => "0010100110000101", 13820 => "1001111011001100", 13821 => "0001101010100000", 13822 => "0001000110001101", 13823 => "1000000011101100", 13824 => "0110111000010001", 13825 => "1011000000011110", 13826 => "1110011001111111", 13827 => "0100011011111100", 13828 => "1101001000111010", 13829 => "0110010010011010", 13830 => "0111011000111010", 13831 => "0100011111110010", 13832 => "1110111000100100", 13833 => "1001100111011111", 13834 => "0110110110110111", 13835 => "1001101111010101", 13836 => "0111110111001001", 13837 => "1100111001010100", 13838 => "1000011001101101", 13839 => "1101111000111111", 13840 => "1000011100101011", 13841 => "0000010010110100", 13842 => "0001101110101100", 13843 => "1101110110111000", 13844 => "0100010000111110", 13845 => "1011100000010001", 13846 => "0010011101101101", 13847 => "0010010110100110", 13848 => "0000110101000111", 13849 => "0111010110110000", 13850 => "1000110111111101", 13851 => "0001100110101010", 13852 => "1011100011011011", 13853 => "1000010011111000", 13854 => "0010010111100111", 13855 => "1001010100001111", 13856 => "0111000010001000", 13857 => "1111110101001110", 13858 => "0010101111111101", 13859 => "0010111011100111", 13860 => "1110011010101100", 13861 => "0100100100101101", 13862 => "0011101010110001", 13863 => "0011000101001111", 13864 => "1000101011111011", 13865 => "0001001011111011", 13866 => "1100011000111111", 13867 => "0111000011000000", 13868 => "0111101000100000", 13869 => "0100110010011110", 13870 => "0111011111111111", 13871 => "1100101111101011", 13872 => "0110100100000101", 13873 => "0100111110101001", 13874 => "1010001100110000", 13875 => "1100111100110101", 13876 => "1000100001111100", 13877 => "1101001010010000", 13878 => "0001011000110100", 13879 => "1111111001001000", 13880 => "1010001101011000", 13881 => "0001011001001011", 13882 => "0010010010110001", 13883 => "0011100011001101", 13884 => "0100001001000001", 13885 => "0101000011001010", 13886 => "0111010110111111", 13887 => "1100101111101011", 13888 => "1010110010010001", 13889 => "0111000010110111", 13890 => "0110101100011011", 13891 => "1000100101011001", 13892 => "1000100011100000", 13893 => "1001011101101110", 13894 => "0100110110011000", 13895 => "1000010111101011", 13896 => "1011000111001010", 13897 => "0111000001010001", 13898 => "1101010110011110", 13899 => "1110010101111001", 13900 => "0010011000110101", 13901 => "0000011100001111", 13902 => "0011001010111100", 13903 => "1100011110011111", 13904 => "0111100101111010", 13905 => "1011101101010110", 13906 => "0100010100111000", 13907 => "1111101011000000", 13908 => "0010110100101101", 13909 => "0101100000000010", 13910 => "1110011010001100", 13911 => "1010010101001110", 13912 => "0111111000011101", 13913 => "0000010001011111", 13914 => "1101011101110110", 13915 => "0111011001011101", 13916 => "1010110001001101", 13917 => "1010100011011000", 13918 => "1011110110010110", 13919 => "0010000100110011", 13920 => "1011011100001000", 13921 => "1001101001001101", 13922 => "0110100111111000", 13923 => "1000010110111111", 13924 => "1000111111100001", 13925 => "1111100100101000", 13926 => "1111111011101000", 13927 => "0111110000010101", 13928 => "1101001111011011", 13929 => "0101001101000011", 13930 => "0011100110101101", 13931 => "1101001001001100", 13932 => "0100101001010001", 13933 => "1100000000010100", 13934 => "1010000100010101", 13935 => "0100111001000111", 13936 => "0000010110000000", 13937 => "0110010010110101", 13938 => "0000001011101001", 13939 => "1010011000001011", 13940 => "1110011000011010", 13941 => "1000100111000001", 13942 => "1101010100111101", 13943 => "0011000010101110", 13944 => "0011011110101000", 13945 => "0101101010100010", 13946 => "0011011111101000", 13947 => "0011001000001100", 13948 => "0111100011000011", 13949 => "1101100010011111", 13950 => "1111000010010111", 13951 => "1100110110100100", 13952 => "0100110001100000", 13953 => "1000111011010011", 13954 => "0101011101111011", 13955 => "1011010011101011", 13956 => "1111010101110101", 13957 => "1111001000010010", 13958 => "1010011100100011", 13959 => "1101001110101100", 13960 => "1111010010000011", 13961 => "1110011001011101", 13962 => "0001011101110101", 13963 => "1010101111001100", 13964 => "0101011100101001", 13965 => "0011100000000111", 13966 => "1110101111000011", 13967 => "0001110000101111", 13968 => "0110100010110001", 13969 => "1001000010100001", 13970 => "1001100000001010", 13971 => "1111010100010110", 13972 => "0001001111111010", 13973 => "0101110001011111", 13974 => "0001110100101001", 13975 => "0000111101010110", 13976 => "1011011011011101", 13977 => "1001010100010010", 13978 => "1010111101100101", 13979 => "1101000010100100", 13980 => "0011111001000110", 13981 => "1010011101001010", 13982 => "0011111000001001", 13983 => "0000111000000010", 13984 => "0001011110011001", 13985 => "1100010001110010", 13986 => "0011110110011110", 13987 => "1111111001111111", 13988 => "1010000011111001", 13989 => "1100111000011101", 13990 => "1000010000010010", 13991 => "1100001010110010", 13992 => "0110111010001110", 13993 => "1111100000110100", 13994 => "0000001110001110", 13995 => "1100110010110110", 13996 => "0100010001101000", 13997 => "0010000001111101", 13998 => "1100000101110111", 13999 => "1111001110001010", 14000 => "0110000101111011", 14001 => "1100101101000000", 14002 => "1111110110100001", 14003 => "0010101100111001", 14004 => "1010110110100101", 14005 => "0110011001110111", 14006 => "1111100100110101", 14007 => "1001111001000010", 14008 => "0100101101011001", 14009 => "1100001010011111", 14010 => "1011001100011011", 14011 => "0110111000010000", 14012 => "1110110111110011", 14013 => "1000010011001000", 14014 => "0100000101010011", 14015 => "1100100111110010", 14016 => "1101000011011111", 14017 => "1110110101000101", 14018 => "0011100111011000", 14019 => "1100100011100000", 14020 => "1001110001110111", 14021 => "1011000101001001", 14022 => "0010010110000000", 14023 => "0111001110001011", 14024 => "0101010111101011", 14025 => "1101100010111001", 14026 => "0000011110000010", 14027 => "1100001111111111", 14028 => "0100001110111001", 14029 => "1100001100110010", 14030 => "1001010000111101", 14031 => "1000100101000111", 14032 => "0011110000011010", 14033 => "0110100111101010", 14034 => "1111001110010011", 14035 => "0000010101011100", 14036 => "1111000111110100", 14037 => "0110111111101110", 14038 => "1000011100011111", 14039 => "1100101100000100", 14040 => "0011100011111111", 14041 => "0101100100010110", 14042 => "0000000101000010", 14043 => "0001010000000100", 14044 => "1000000100000111", 14045 => "0111000101001110", 14046 => "0011011000100111", 14047 => "1100001110101100", 14048 => "0110111101101101", 14049 => "1001010010010101", 14050 => "1110111110010101", 14051 => "0001101100100101", 14052 => "1110101010100110", 14053 => "0101001011111111", 14054 => "1100010011110100", 14055 => "0000101101110000", 14056 => "0110100011100100", 14057 => "0000111010100110", 14058 => "1000000010001110", 14059 => "1110111011110000", 14060 => "0100000001010100", 14061 => "1101000110110101", 14062 => "0010000110110011", 14063 => "1100110111001101", 14064 => "0001111001011111", 14065 => "1100110110000001", 14066 => "1110010001100001", 14067 => "1101001000100010", 14068 => "0010100101011001", 14069 => "1001000000100110", 14070 => "1001010110001011", 14071 => "1100001001011101", 14072 => "0111110111100000", 14073 => "0001001110000110", 14074 => "0110101100001001", 14075 => "1000011111001110", 14076 => "0110000111111010", 14077 => "1111100010110010", 14078 => "0000011110010110", 14079 => "1000010011001100", 14080 => "1011101000100110", 14081 => "0001100100001101", 14082 => "1110100110010101", 14083 => "0111001001000100", 14084 => "1111000100101011", 14085 => "0011110111110101", 14086 => "1000000000010001", 14087 => "1001010100111010", 14088 => "1011110001001100", 14089 => "1010100000111000", 14090 => "1010001100011110", 14091 => "1101100001111000", 14092 => "1010000110000111", 14093 => "1111100101110010", 14094 => "1101011110110100", 14095 => "0011111111010101", 14096 => "0101010010110101", 14097 => "1001110011100011", 14098 => "1111000011101111", 14099 => "0101101110101101", 14100 => "0100010111000000", 14101 => "1100110100111011", 14102 => "1110111011010000", 14103 => "0101000101011110", 14104 => "0001010111110100", 14105 => "0111110000000110", 14106 => "1101100111100001", 14107 => "1111111101100000", 14108 => "0110101001111100", 14109 => "0010101010000000", 14110 => "1000101011011001", 14111 => "1011101101010010", 14112 => "1111000100011011", 14113 => "1000101010010011", 14114 => "0110100101110100", 14115 => "1000001101011100", 14116 => "0000001101111111", 14117 => "1011110100001111", 14118 => "0011000011000110", 14119 => "0000011001101000", 14120 => "0111100000001110", 14121 => "1110001100111011", 14122 => "1101000111101101", 14123 => "1101010111110111", 14124 => "0110100011100110", 14125 => "1111000101101101", 14126 => "0011011010101101", 14127 => "1111010010010000", 14128 => "0001110100100010", 14129 => "0011100110011100", 14130 => "0101000000011000", 14131 => "0111110101011111", 14132 => "1011101101111000", 14133 => "1101001011110011", 14134 => "0000000111011010", 14135 => "1100010100101110", 14136 => "1001110000110100", 14137 => "1110011101110001", 14138 => "0001001110110001", 14139 => "1111010100111011", 14140 => "0111111100100010", 14141 => "1000000110001000", 14142 => "1110011110110110", 14143 => "1101101110011111", 14144 => "0001111011011000", 14145 => "1101010000100110", 14146 => "0011000110010001", 14147 => "1011101100101001", 14148 => "1011010000101110", 14149 => "0000000111111011", 14150 => "1100111100111010", 14151 => "0111110111001110", 14152 => "0010101011010111", 14153 => "1010000000101101", 14154 => "0001100100111001", 14155 => "0110111000011110", 14156 => "0100000100001011", 14157 => "0110100001110010", 14158 => "1001101001001111", 14159 => "1000111110110010", 14160 => "0011111111100010", 14161 => "1011001010000100", 14162 => "1000011000011011", 14163 => "1000110101100100", 14164 => "1010010001101010", 14165 => "0101110100111001", 14166 => "1111010010000010", 14167 => "0110101100110110", 14168 => "0100010100010001", 14169 => "1101000010001000", 14170 => "0100100111111011", 14171 => "1111000011100110", 14172 => "0101110111011011", 14173 => "1001010000111101", 14174 => "1100100110011011", 14175 => "0000110011110100", 14176 => "1100101101011011", 14177 => "0100100110110101", 14178 => "0000101111000000", 14179 => "1100111010100001", 14180 => "0011001000010000", 14181 => "1101100100111111", 14182 => "0001101000101100", 14183 => "1000111011111000", 14184 => "1101101100000000", 14185 => "0000000110110001", 14186 => "0101000000000011", 14187 => "1011001010101100", 14188 => "0100101000110111", 14189 => "1010101011101000", 14190 => "0110000101011100", 14191 => "0100111000001110", 14192 => "1000000000011011", 14193 => "1000101001101010", 14194 => "0110100100010101", 14195 => "0000000110100110", 14196 => "0001101101111100", 14197 => "1010101000111001", 14198 => "1111110011010110", 14199 => "0001000111011010", 14200 => "1111011100100111", 14201 => "0011010010100110", 14202 => "0011000001101000", 14203 => "1110101100001011", 14204 => "1011000010010100", 14205 => "1100111100011000", 14206 => "0100100000100111", 14207 => "0000001011010010", 14208 => "1111000101110101", 14209 => "1000111110100110", 14210 => "1001100101001011", 14211 => "0001001110110110", 14212 => "1010011001000001", 14213 => "0110010111101001", 14214 => "1010011100000010", 14215 => "0111011010111110", 14216 => "1010111100101101", 14217 => "0010001101011010", 14218 => "0001011010101110", 14219 => "1111111000101011", 14220 => "1100011110001001", 14221 => "1111100111111000", 14222 => "1011011011100011", 14223 => "1001101001100000", 14224 => "1101011111011111", 14225 => "0110000011110101", 14226 => "0111111000101101", 14227 => "1111101110000001", 14228 => "0111100111011000", 14229 => "0111111001001101", 14230 => "0001000110100100", 14231 => "1111000010100011", 14232 => "1110000011100100", 14233 => "1111001000001010", 14234 => "0110011011100001", 14235 => "1111111010111010", 14236 => "1011010110011010", 14237 => "1010001110000011", 14238 => "1101000100001110", 14239 => "1100110111011001", 14240 => "1000011001101101", 14241 => "0000011110000100", 14242 => "1100101101001101", 14243 => "0111110111101001", 14244 => "1100100110100111", 14245 => "1010000011001001", 14246 => "0111100001000000", 14247 => "1000100000011110", 14248 => "1011001010001000", 14249 => "1000111001100100", 14250 => "1100000010001001", 14251 => "0000001000100000", 14252 => "0000101110001001", 14253 => "1010100110110110", 14254 => "1101010000100101", 14255 => "1111111001101101", 14256 => "0111101011110101", 14257 => "1011011010100100", 14258 => "1000010000111000", 14259 => "1100001011011111", 14260 => "0001001001110001", 14261 => "1010101111110011", 14262 => "0101001111001011", 14263 => "1111001011000001", 14264 => "0110101001000111", 14265 => "1100010000100001", 14266 => "0001010000101001", 14267 => "1100101001101001", 14268 => "1011011001001011", 14269 => "0101010011011101", 14270 => "0011010001100010", 14271 => "1001000010000001", 14272 => "1001110101011001", 14273 => "1101100110001100", 14274 => "1110000000101110", 14275 => "1000001111111011", 14276 => "0011111101001111", 14277 => "0101001010000010", 14278 => "0110111101010111", 14279 => "1000001010110000", 14280 => "0101110100111001", 14281 => "0001110101001101", 14282 => "1100101100010101", 14283 => "0101000011010011", 14284 => "1001101111011011", 14285 => "1101010010001110", 14286 => "1110101001100011", 14287 => "1010001111010001", 14288 => "0101100100000111", 14289 => "0101001101000100", 14290 => "1101100000011111", 14291 => "0101111010001111", 14292 => "1110010011100010", 14293 => "1110001011000011", 14294 => "1100110111000111", 14295 => "1101000010000001", 14296 => "1011001001010111", 14297 => "0111000111100100", 14298 => "1110011101111000", 14299 => "1111111010000011", 14300 => "0100010111111110", 14301 => "1010011000001101", 14302 => "1000110101001010", 14303 => "0011001111001101", 14304 => "0011011100100100", 14305 => "1110000011011011", 14306 => "1001010100010011", 14307 => "1010101110110110", 14308 => "1110111001011111", 14309 => "1111011010101000", 14310 => "1100101110000000", 14311 => "0100010111101100", 14312 => "0010011010001011", 14313 => "0111011011011001", 14314 => "0100011100011110", 14315 => "1111001111101000", 14316 => "0010010100110011", 14317 => "1001001100011100", 14318 => "0100000100110000", 14319 => "0010110101110011", 14320 => "1001010001100010", 14321 => "1101001100100101", 14322 => "1000011011111111", 14323 => "1010110011110101", 14324 => "1011011110011000", 14325 => "0100011110110110", 14326 => "0111010000001011", 14327 => "1000010100100000", 14328 => "0010111100001110", 14329 => "0000110000001110", 14330 => "1111001100011100", 14331 => "0011100100010110", 14332 => "0011010000110010", 14333 => "0010101011010010", 14334 => "0011010100100111", 14335 => "0101100111010100", 14336 => "0100010101001101", 14337 => "0001111001101110", 14338 => "0111100001011010", 14339 => "0000101100010101", 14340 => "1000110011011001", 14341 => "0100010100101101", 14342 => "0110010011010101", 14343 => "1000010011000110", 14344 => "1101011000001000", 14345 => "1010110000110010", 14346 => "0110001000111000", 14347 => "1111001110110100", 14348 => "0010000100101010", 14349 => "0010010101111101", 14350 => "0100101001011100", 14351 => "0000101010000010", 14352 => "0010010000001111", 14353 => "0011101010001100", 14354 => "0010001100101100", 14355 => "0000010011100111", 14356 => "1001111110101001", 14357 => "0000000111000111", 14358 => "1001111011000011", 14359 => "1110000101000010", 14360 => "1000101001110000", 14361 => "1111101001100111", 14362 => "1001101010000001", 14363 => "1000101101011011", 14364 => "0110010111001101", 14365 => "1111100001001111", 14366 => "0111100111101000", 14367 => "0110110100110001", 14368 => "1100001100011011", 14369 => "0010001110001111", 14370 => "0101001000101011", 14371 => "0000101000010101", 14372 => "1010110000000101", 14373 => "0100000000011111", 14374 => "1000010010010101", 14375 => "0011100001010111", 14376 => "0000011100001000", 14377 => "1100100001101110", 14378 => "1110111000111000", 14379 => "1000100101011010", 14380 => "0001010110010011", 14381 => "0010001011111100", 14382 => "1111101100100001", 14383 => "1011011101000111", 14384 => "0001111001100010", 14385 => "1010010000110111", 14386 => "0101000001001111", 14387 => "1100100001010111", 14388 => "1111111100100010", 14389 => "0010001010000101", 14390 => "1011000010010100", 14391 => "1010100001001111", 14392 => "1000011100101110", 14393 => "0001000100010100", 14394 => "1111100010110101", 14395 => "0011010011000111", 14396 => "0111100010100010", 14397 => "1001010001011101", 14398 => "1010000110101110", 14399 => "1001001110010000", 14400 => "1100101100000101", 14401 => "1001000010001110", 14402 => "1000001111001110", 14403 => "0100111011100110", 14404 => "1011000010001000", 14405 => "1111011101111101", 14406 => "0010100100010000", 14407 => "0001011001111001", 14408 => "1001100000110100", 14409 => "1111110111011101", 14410 => "1011111111000100", 14411 => "1100001111010110", 14412 => "1011100001110001", 14413 => "1110111001100100", 14414 => "0010101011100010", 14415 => "0110000000111111", 14416 => "0101110001011010", 14417 => "1000010011101100", 14418 => "1001111100010111", 14419 => "1110111101011100", 14420 => "0101100010011110", 14421 => "0010011010001100", 14422 => "0010100110010011", 14423 => "1100011010100000", 14424 => "1010011110111001", 14425 => "1001101000010011", 14426 => "0000110111110000", 14427 => "1011111101111101", 14428 => "1000110011111100", 14429 => "1001101000111000", 14430 => "1000010110000100", 14431 => "1101000000011001", 14432 => "0011100110110010", 14433 => "1000010110100111", 14434 => "0110111001001010", 14435 => "0000111101100010", 14436 => "1100000010000010", 14437 => "1010001000110001", 14438 => "0110100111111100", 14439 => "0100010000110111", 14440 => "0100110100001110", 14441 => "0000010100100010", 14442 => "1010011000010101", 14443 => "1111111101000111", 14444 => "0001010101110011", 14445 => "0001001100011110", 14446 => "0011100011111000", 14447 => "0100111100011101", 14448 => "0111101101100011", 14449 => "1111010101111100", 14450 => "1000110110101000", 14451 => "1001011111000110", 14452 => "1001000100001001", 14453 => "0110011010000110", 14454 => "1101111001001111", 14455 => "1101000100011001", 14456 => "1101100111101100", 14457 => "1111101111110000", 14458 => "0110100110110001", 14459 => "0101111001001110", 14460 => "0100000010101101", 14461 => "1011000111101010", 14462 => "1001100101001011", 14463 => "0010011010101000", 14464 => "0111001000000000", 14465 => "1001101011000010", 14466 => "0111001011111010", 14467 => "0110001101111011", 14468 => "0101000000101100", 14469 => "0100001011001001", 14470 => "0111010010111001", 14471 => "0000111100100011", 14472 => "1111110111011111", 14473 => "1110010111111111", 14474 => "1100000001101010", 14475 => "1000110001001111", 14476 => "0100101101010001", 14477 => "0011001000100011", 14478 => "1010101110111111", 14479 => "0000000111000111", 14480 => "1110100011000011", 14481 => "1100100100010000", 14482 => "1000111111011111", 14483 => "0111101100001011", 14484 => "1100101111010111", 14485 => "1011111100100001", 14486 => "0111110110111001", 14487 => "0010000101001111", 14488 => "1100100111000011", 14489 => "1010100000011011", 14490 => "0000011101111001", 14491 => "0001111010000110", 14492 => "1111001100000110", 14493 => "0011110000010100", 14494 => "1111010101001110", 14495 => "0100101011101001", 14496 => "1110101101001111", 14497 => "1010111101011010", 14498 => "0101000001110000", 14499 => "1011010100110110", 14500 => "1101101100001100", 14501 => "1010110011011011", 14502 => "1011100010100011", 14503 => "1101100010001010", 14504 => "0111111000110101", 14505 => "1111110110111011", 14506 => "0111100000110111", 14507 => "1010000010010101", 14508 => "0010000100100000", 14509 => "0000011001101101", 14510 => "1100011101100010", 14511 => "1000010011011010", 14512 => "1101001001111011", 14513 => "1011011011100101", 14514 => "1101000001110101", 14515 => "1000111000101101", 14516 => "1001010110000101", 14517 => "1101011110111110", 14518 => "0101111000111010", 14519 => "1011110110001011", 14520 => "1110110110110001", 14521 => "1001100101111111", 14522 => "0011001001101011", 14523 => "1111011011101011", 14524 => "1111100110001110", 14525 => "0101011001110111", 14526 => "1010001001100000", 14527 => "1110110111011010", 14528 => "1010100000111000", 14529 => "0000010001100000", 14530 => "0111011101110110", 14531 => "1100100101001011", 14532 => "0101101011101101", 14533 => "1110010010011000", 14534 => "1000010110100110", 14535 => "1101001011101111", 14536 => "1000101101001110", 14537 => "1110100011101111", 14538 => "1011000111011010", 14539 => "1001000110011100", 14540 => "0101100001111111", 14541 => "0000010100000011", 14542 => "1100001101001100", 14543 => "1010101100010100", 14544 => "0101001111111001", 14545 => "0000011110110111", 14546 => "1010010011000101", 14547 => "0111010110000100", 14548 => "1101001100101100", 14549 => "1010000100001000", 14550 => "1101011111010110", 14551 => "0001111000011000", 14552 => "0010110001101110", 14553 => "0110010100101111", 14554 => "0010001110010011", 14555 => "0100010001010000", 14556 => "1000010100001011", 14557 => "0010100111111100", 14558 => "0010010111110001", 14559 => "1110010010101010", 14560 => "0110000011001101", 14561 => "1101010111000110", 14562 => "0011101010010011", 14563 => "0110110001010000", 14564 => "0110011110001101", 14565 => "0001000011100001", 14566 => "0010101001100001", 14567 => "1111000101100101", 14568 => "0011000101011000", 14569 => "1101001010101000", 14570 => "0000111110101100", 14571 => "1000110100100000", 14572 => "1101111111101111", 14573 => "0110100000010110", 14574 => "0000110110100101", 14575 => "1001010111000010", 14576 => "0101011001011111", 14577 => "0010001110001011", 14578 => "0110011001010010", 14579 => "1000010011011111", 14580 => "0110111011001100", 14581 => "1111001101100010", 14582 => "0011010110111101", 14583 => "1100001010011100", 14584 => "0111101011011011", 14585 => "1111001110110001", 14586 => "1010111011111000", 14587 => "1011010100111111", 14588 => "0010100011001010", 14589 => "1010000100101010", 14590 => "1000011111001111", 14591 => "1000000001010100", 14592 => "1110000110111010", 14593 => "0011111010011110", 14594 => "0011101111001111", 14595 => "1000000011010011", 14596 => "1010100111111000", 14597 => "0010000001001111", 14598 => "1010101110111010", 14599 => "0111111110010011", 14600 => "1100111100011001", 14601 => "0111100111111010", 14602 => "0000101001011110", 14603 => "0000111100001010", 14604 => "0000000011110001", 14605 => "1100100100111110", 14606 => "1011101010101101", 14607 => "0010101101111110", 14608 => "1001101110000011", 14609 => "1010000110001100", 14610 => "1000000101000001", 14611 => "0111011001101001", 14612 => "0100101010000010", 14613 => "0101110100110110", 14614 => "0100111110011111", 14615 => "0111001000110101", 14616 => "0010011101111110", 14617 => "0101011110100101", 14618 => "0100111101101000", 14619 => "1011011001100100", 14620 => "1000100111000110", 14621 => "0100100010110010", 14622 => "1000100100010101", 14623 => "1011011101111010", 14624 => "0111111100011001", 14625 => "0100101111110011", 14626 => "1011101110100101", 14627 => "1001011101101100", 14628 => "0000010011100111", 14629 => "1111000111010110", 14630 => "1110110110011011", 14631 => "1110000110110011", 14632 => "1010111011010111", 14633 => "0000110100000100", 14634 => "1010101111010100", 14635 => "0101100000010101", 14636 => "0001000110100010", 14637 => "0011010111011010", 14638 => "0000011100001100", 14639 => "0001101100001111", 14640 => "0111010100000100", 14641 => "1000000011010010", 14642 => "1110101110111110", 14643 => "1100010110111100", 14644 => "1001001001010010", 14645 => "1101110101000001", 14646 => "0110110000000100", 14647 => "1010000001000111", 14648 => "0010101011001100", 14649 => "0011101011110111", 14650 => "1001111111110110", 14651 => "1000110001110111", 14652 => "0101001001101110", 14653 => "0010110000001010", 14654 => "0110000010101000", 14655 => "0110110011100111", 14656 => "0000011011111000", 14657 => "0001010010011100", 14658 => "0111011111101110", 14659 => "1110001111101010", 14660 => "1100101010011011", 14661 => "1010110010111011", 14662 => "1101001100110110", 14663 => "1110100010100000", 14664 => "0101100001010001", 14665 => "0011110100110100", 14666 => "0001111001000110", 14667 => "0100011110110011", 14668 => "1011011001101101", 14669 => "0111111110001000", 14670 => "0110000011010100", 14671 => "1101100011000011", 14672 => "0100100011110111", 14673 => "0101010000101111", 14674 => "0000110100001010", 14675 => "0110101000001100", 14676 => "0100000000111011", 14677 => "1010110101100010", 14678 => "0110111111111110", 14679 => "0101000010011001", 14680 => "0100011100001110", 14681 => "0101001100011010", 14682 => "0011010000110101", 14683 => "1100000010100111", 14684 => "1001111110100100", 14685 => "1011001011101111", 14686 => "0100111101110100", 14687 => "0101101011100011", 14688 => "1100000011100001", 14689 => "1101010000001100", 14690 => "1110001011101110", 14691 => "0100101000111110", 14692 => "0001010001111010", 14693 => "1101000011000110", 14694 => "0111001100001110", 14695 => "0000000000000000", 14696 => "1101011000011101", 14697 => "0100000010111000", 14698 => "1101011001100110", 14699 => "1011000010100001", 14700 => "0000000100010101", 14701 => "0101110101000110", 14702 => "1110010110100101", 14703 => "1101100111001110", 14704 => "0101000010100001", 14705 => "1001110110011101", 14706 => "0001111010011111", 14707 => "0011101011101011", 14708 => "0101001101101101", 14709 => "1111010000001111", 14710 => "0000100001010011", 14711 => "0111011111011011", 14712 => "1100111111101010", 14713 => "1111010010100011", 14714 => "1110011011111100", 14715 => "0001101110001100", 14716 => "1001001100101011", 14717 => "0111111011111110", 14718 => "0010101000011100", 14719 => "0111010010011010", 14720 => "1110110001001001", 14721 => "0000111101101100", 14722 => "1010101001111110", 14723 => "1100001011010011", 14724 => "1001001011001000", 14725 => "1101110000001101", 14726 => "0100101110111001", 14727 => "0101001110000010", 14728 => "1011001101111000", 14729 => "1011100001001000", 14730 => "0011110110010100", 14731 => "0010100111101011", 14732 => "1010011100100011", 14733 => "1111101110011110", 14734 => "0011101100001010", 14735 => "0000110011010010", 14736 => "1101100000000101", 14737 => "1100001111010111", 14738 => "0001100100001010", 14739 => "1010111010010110", 14740 => "1101001000011101", 14741 => "0111001111000101", 14742 => "0111101111000101", 14743 => "0010001011000110", 14744 => "0100011011100010", 14745 => "1111011001011110", 14746 => "1000101000100011", 14747 => "1110010010100011", 14748 => "1110101000001101", 14749 => "0011101101001010", 14750 => "0100111110000010", 14751 => "1010100110101010", 14752 => "1101010010000100", 14753 => "1111111000110001", 14754 => "1100101001100010", 14755 => "1101101110010101", 14756 => "0010101001011000", 14757 => "1110001101011011", 14758 => "0101001010010101", 14759 => "0110011110010000", 14760 => "1110110101110000", 14761 => "0110001110110110", 14762 => "1111110000011000", 14763 => "1001001000011011", 14764 => "1110110001110010", 14765 => "0111010011100010", 14766 => "1011000100011111", 14767 => "0110011000001011", 14768 => "0110101001110001", 14769 => "0100010100101100", 14770 => "1111000100111100", 14771 => "0000000111111100", 14772 => "1000000111111110", 14773 => "0101111011110100", 14774 => "1111001010100101", 14775 => "0111100101100101", 14776 => "0011011001000001", 14777 => "1101011101111110", 14778 => "0000110000101001", 14779 => "0011100010111101", 14780 => "0111000001011110", 14781 => "1101111011101010", 14782 => "0111001001101000", 14783 => "0000001101000001", 14784 => "1100001100001111", 14785 => "0111010000001000", 14786 => "0110010010100011", 14787 => "0110001001001001", 14788 => "0001010101110111", 14789 => "0001101001011110", 14790 => "0101111101001001", 14791 => "0100101110001110", 14792 => "0110000000010100", 14793 => "0000110100000000", 14794 => "0001001011000111", 14795 => "0001101100100011", 14796 => "1011001011000111", 14797 => "1011100100011001", 14798 => "0000111110110100", 14799 => "1100001101011001", 14800 => "1001011111000000", 14801 => "0111001110011010", 14802 => "1001000101010010", 14803 => "0111000100001110", 14804 => "1011011001110101", 14805 => "1010110000111101", 14806 => "0111010111001001", 14807 => "1101110010000001", 14808 => "1000010110011111", 14809 => "1111101110011110", 14810 => "0010111010000100", 14811 => "1010101001110000", 14812 => "1111100010110100", 14813 => "1001100100010111", 14814 => "0010000111101000", 14815 => "1011101011100110", 14816 => "1110011100101100", 14817 => "1111111011011110", 14818 => "1110011011001011", 14819 => "1101001101011110", 14820 => "1011000001110100", 14821 => "0100110111000001", 14822 => "0111111001111110", 14823 => "0011000111011100", 14824 => "0011001000100100", 14825 => "0110011000011000", 14826 => "1010101001001001", 14827 => "0110101011000111", 14828 => "0100011010010011", 14829 => "1000100111100111", 14830 => "1000010100000111", 14831 => "0101101011001111", 14832 => "0100010111000010", 14833 => "1100110010011001", 14834 => "0111010000100011", 14835 => "0000111011000110", 14836 => "1000001110011111", 14837 => "1111100011011001", 14838 => "1001000001110110", 14839 => "0101000101100000", 14840 => "1101101101111110", 14841 => "1111011010111110", 14842 => "0000011000000100", 14843 => "0001101100101111", 14844 => "1011101001001010", 14845 => "1011011000100111", 14846 => "0010010000010000", 14847 => "1111000110000000", 14848 => "1101100110100111", 14849 => "1100110110001101", 14850 => "0100111111110000", 14851 => "0001000001101001", 14852 => "0101011001100101", 14853 => "0111000001100001", 14854 => "1010000000010001", 14855 => "1111100011101110", 14856 => "0101110010000011", 14857 => "1000000010110111", 14858 => "1000011010101000", 14859 => "1010110111010011", 14860 => "1001110111111001", 14861 => "1000110100100100", 14862 => "0111000010110111", 14863 => "1010001011000100", 14864 => "1100010101001011", 14865 => "0101010110111000", 14866 => "0010100010010101", 14867 => "1010011101011010", 14868 => "1011010010001110", 14869 => "1000101001001011", 14870 => "0001011110011110", 14871 => "1000101110010010", 14872 => "1110001000000110", 14873 => "1100001111111001", 14874 => "0101100000100001", 14875 => "0001111110101110", 14876 => "1111100110101001", 14877 => "0001001010011100", 14878 => "1011110100011110", 14879 => "0101101111001101", 14880 => "0110100011010010", 14881 => "1101001100011111", 14882 => "1011010001101100", 14883 => "0010110011011100", 14884 => "1110110011100110", 14885 => "1110010010000011", 14886 => "1100100110101100", 14887 => "0000100010011111", 14888 => "0111101100110110", 14889 => "1110000101110001", 14890 => "0111010101010111", 14891 => "0101110011001100", 14892 => "0010001010011010", 14893 => "0100110101111011", 14894 => "1001111011110001", 14895 => "0000000111000010", 14896 => "1000001011101001", 14897 => "0100000100110111", 14898 => "0111111010111000", 14899 => "1011000010001100", 14900 => "1101001100001111", 14901 => "1110011110001111", 14902 => "1000100100100100", 14903 => "0010111011110111", 14904 => "1100010010100110", 14905 => "1101110100101100", 14906 => "0011010011000011", 14907 => "1000000001101111", 14908 => "0001011110011000", 14909 => "1111110001101100", 14910 => "0000100110111010", 14911 => "0011010001101100", 14912 => "1010110010011001", 14913 => "0110111100100110", 14914 => "0111110001100110", 14915 => "0100011001010101", 14916 => "1111111010000001", 14917 => "1001001100011001", 14918 => "1101010111101000", 14919 => "0000000100011111", 14920 => "0111010000010101", 14921 => "0101101000010100", 14922 => "1100111010010100", 14923 => "0011011001010010", 14924 => "1101011000111111", 14925 => "0110110100010111", 14926 => "0010001001101010", 14927 => "0000101010111101", 14928 => "0010001101100110", 14929 => "0011111101101010", 14930 => "0110011101111100", 14931 => "0100100100001010", 14932 => "0111010001011110", 14933 => "0101111000011001", 14934 => "0110100100101000", 14935 => "1011001111000000", 14936 => "0001111101100011", 14937 => "1001111011101100", 14938 => "1010000111111010", 14939 => "1001001010100000", 14940 => "1011110011111001", 14941 => "1001000010011101", 14942 => "0010111110010011", 14943 => "1100000001101101", 14944 => "0111111101101101", 14945 => "0010011011011110", 14946 => "0100111111110000", 14947 => "0001001001101111", 14948 => "1111011001101011", 14949 => "1010011100000110", 14950 => "0010010001110000", 14951 => "1010111000111110", 14952 => "0000000100110011", 14953 => "0111110011001101", 14954 => "0100111001101100", 14955 => "0001001001101010", 14956 => "0000001000011100", 14957 => "0001111101010010", 14958 => "0001001101111000", 14959 => "0110011011100010", 14960 => "1000110001110000", 14961 => "0000111011111000", 14962 => "0011111110101001", 14963 => "1100000101010011", 14964 => "0010011011011001", 14965 => "1011100011111000", 14966 => "0000101001010010", 14967 => "0000010001100101", 14968 => "1010101111111011", 14969 => "1000100100110100", 14970 => "1010111101110111", 14971 => "0011010111101111", 14972 => "1011001111010011", 14973 => "1010111000001001", 14974 => "1011010101111010", 14975 => "0100110011000101", 14976 => "1010111011001010", 14977 => "0100011100101110", 14978 => "1001101010100110", 14979 => "0011011100111110", 14980 => "1110110111000110", 14981 => "0111000101100110", 14982 => "0010100101100101", 14983 => "0111110010000011", 14984 => "1100001010010101", 14985 => "1100011110001001", 14986 => "0010010001000111", 14987 => "0001100101010001", 14988 => "0111010100100001", 14989 => "1101010100110100", 14990 => "1101101000100111", 14991 => "0010101001100001", 14992 => "1000111101100011", 14993 => "1010011000001111", 14994 => "1111111000110001", 14995 => "1011000101100011", 14996 => "0010101111110000", 14997 => "0111011010111110", 14998 => "1110100001100101", 14999 => "1100010000001100", 15000 => "1100100111100011", 15001 => "0110001001100110", 15002 => "1110010001001110", 15003 => "1100101101100100", 15004 => "0000000001101100", 15005 => "1111111010011000", 15006 => "1010011110001011", 15007 => "0011111001111000", 15008 => "1001100101101000", 15009 => "1000000001000010", 15010 => "0110001111001010", 15011 => "0000110100000110", 15012 => "1000011011010001", 15013 => "0001011010001101", 15014 => "0101100011101001", 15015 => "0010010110101001", 15016 => "1000011010101011", 15017 => "0110001100100101", 15018 => "0000001001100010", 15019 => "0111101011110110", 15020 => "1001011101100101", 15021 => "0000010000011000", 15022 => "1001011000100000", 15023 => "1100100011110100", 15024 => "0101110000101101", 15025 => "1110100100101001", 15026 => "1011100010011111", 15027 => "0110100001000011", 15028 => "1111111011001101", 15029 => "1010111111101011", 15030 => "0100101000100110", 15031 => "0111011001010100", 15032 => "0100111110001101", 15033 => "0011011101101101", 15034 => "1010001011100100", 15035 => "0101110101110110", 15036 => "1110001111111010", 15037 => "0000000010000001", 15038 => "1001010111110001", 15039 => "0111011111101100", 15040 => "1010011110100011", 15041 => "0010010010000010", 15042 => "0100101111110110", 15043 => "0100101111100101", 15044 => "0101010011000111", 15045 => "0100010000100101", 15046 => "1110001111011001", 15047 => "0010010111000011", 15048 => "0000011011010100", 15049 => "1100111001100101", 15050 => "1111000000001011", 15051 => "0010001000000111", 15052 => "1011011101000000", 15053 => "1010000010000100", 15054 => "0010111010110110", 15055 => "0000011101011110", 15056 => "0001100000101011", 15057 => "1110111111010111", 15058 => "0011011000101010", 15059 => "0000000011010011", 15060 => "1110011110111101", 15061 => "0011110000010001", 15062 => "1100110110110010", 15063 => "0001101100110110", 15064 => "1111000010101010", 15065 => "0101101001000011", 15066 => "0101000110011111", 15067 => "1100111011101101", 15068 => "1001000010001111", 15069 => "1011100100111001", 15070 => "0010010101101001", 15071 => "0010110000000010", 15072 => "1000101100101011", 15073 => "0000010110011011", 15074 => "1001000001011011", 15075 => "0011100001110111", 15076 => "0010001011000001", 15077 => "1010011000111011", 15078 => "0010010100101101", 15079 => "0011000000000010", 15080 => "1001010111111111", 15081 => "0110111010010100", 15082 => "1111101101111011", 15083 => "1111110100111010", 15084 => "1101010110100001", 15085 => "1011010010110001", 15086 => "0000100010111011", 15087 => "0111101110001000", 15088 => "1010001100000110", 15089 => "0010111000111110", 15090 => "0100101100101101", 15091 => "1100111111011010", 15092 => "0000101010111001", 15093 => "1000001010100111", 15094 => "0110110011000011", 15095 => "1011010000010000", 15096 => "1011001100101111", 15097 => "1110000110001000", 15098 => "0001101101101110", 15099 => "0111110111101110", 15100 => "1001001110010011", 15101 => "1010100110101001", 15102 => "0000010000011110", 15103 => "0101001001101111", 15104 => "1011101111100110", 15105 => "1100111101100000", 15106 => "0111100110001111", 15107 => "0000101101010000", 15108 => "0011110100101111", 15109 => "1010100001110110", 15110 => "0100001000010110", 15111 => "0110110111100010", 15112 => "0001111100010010", 15113 => "1111001011000011", 15114 => "1011101100001101", 15115 => "1110001001011110", 15116 => "1001001111010110", 15117 => "1010001111011010", 15118 => "0100101001010100", 15119 => "0001110010101010", 15120 => "0011110001010010", 15121 => "1011110100110001", 15122 => "0110000000111111", 15123 => "0100010000011111", 15124 => "1001101111001110", 15125 => "0101011010101000", 15126 => "1011100101100110", 15127 => "0001111001100000", 15128 => "1111101100100111", 15129 => "0111011001100100", 15130 => "1010111000000000", 15131 => "1000000111101010", 15132 => "1100111010101001", 15133 => "0001101111110001", 15134 => "1101110011101001", 15135 => "0100111001110110", 15136 => "1101001001001001", 15137 => "1010001110010110", 15138 => "0010100111101111", 15139 => "0101111001011000", 15140 => "1010001101011010", 15141 => "0010010010001111", 15142 => "0110100110101001", 15143 => "0011011100010010", 15144 => "1101010101000010", 15145 => "0000110010110110", 15146 => "1010111001101000", 15147 => "1111100010111100", 15148 => "0000001000110001", 15149 => "1101010110010111", 15150 => "0110010111001110", 15151 => "1101101000110001", 15152 => "1101011111000001", 15153 => "1100110010010100", 15154 => "1101001001001111", 15155 => "0100101101000010", 15156 => "1111011000011101", 15157 => "0101011110110101", 15158 => "1000101000110000", 15159 => "0100100110110010", 15160 => "0011010111111000", 15161 => "1101011010011001", 15162 => "1011101010001101", 15163 => "1101000000111111", 15164 => "1111101100010111", 15165 => "1101111110010110", 15166 => "0100110100100111", 15167 => "0010111111110101", 15168 => "0111100011000110", 15169 => "1101111011101011", 15170 => "1100001011111111", 15171 => "1101001010100110", 15172 => "0011110001110001", 15173 => "1100100101110010", 15174 => "0100111001010000", 15175 => "1011101011011110", 15176 => "1110100111110101", 15177 => "0001010100110111", 15178 => "0000110011110000", 15179 => "0111001110000011", 15180 => "0111011101111110", 15181 => "0100111011011011", 15182 => "1011001101110101", 15183 => "1000100000100101", 15184 => "1001011001011001", 15185 => "1110011001101000", 15186 => "0010011110110111", 15187 => "1100001000010010", 15188 => "1001011010001001", 15189 => "0011110010001001", 15190 => "0101111000000010", 15191 => "0110101001011100", 15192 => "1001110101110110", 15193 => "1100101101111100", 15194 => "1111001110100011", 15195 => "1111110001110101", 15196 => "0110111010100101", 15197 => "1101110011111110", 15198 => "0000111101000110", 15199 => "0010011011010010", 15200 => "0010101011101011", 15201 => "0010111101000110", 15202 => "0010001111001111", 15203 => "0100101010011111", 15204 => "1101001110101011", 15205 => "1001000000111110", 15206 => "1000011111100100", 15207 => "0101011001111101", 15208 => "0100111111111010", 15209 => "0000100001001110", 15210 => "0110100100110010", 15211 => "1011000000010101", 15212 => "0100010111011111", 15213 => "1010011010010011", 15214 => "1111010001011100", 15215 => "1000000011111011", 15216 => "0101001111101010", 15217 => "1110111101110100", 15218 => "1101011101100000", 15219 => "0100101100001100", 15220 => "0001110000100010", 15221 => "1110011101101011", 15222 => "0010001110001101", 15223 => "0010110001110101", 15224 => "1011010010111100", 15225 => "1111111001110011", 15226 => "1000101001100001", 15227 => "0011111000111000", 15228 => "0010001111101000", 15229 => "1111010100001011", 15230 => "1011001100000011", 15231 => "0111100111011101", 15232 => "0111111011010110", 15233 => "0111111011011111", 15234 => "1000000101111111", 15235 => "0000000010010111", 15236 => "0101000011110100", 15237 => "1011011110001100", 15238 => "0111011010000111", 15239 => "1011001111001111", 15240 => "1110000010010110", 15241 => "1110001011100001", 15242 => "0011000000111111", 15243 => "1110011110000011", 15244 => "1110111010111100", 15245 => "1001011110101111", 15246 => "0100111110000101", 15247 => "1011110011000100", 15248 => "1010100000011001", 15249 => "0100101001110111", 15250 => "1011010000111110", 15251 => "1101011111101010", 15252 => "0101111011101110", 15253 => "1111101110111110", 15254 => "0010100011010110", 15255 => "0001111111100110", 15256 => "1011010010010111", 15257 => "0111010011111011", 15258 => "0110110100011000", 15259 => "0100100000001101", 15260 => "0100110001010101", 15261 => "1101001001111010", 15262 => "0000111111101001", 15263 => "1000101011010000", 15264 => "1011100001100011", 15265 => "0100001101111010", 15266 => "0000000001111100", 15267 => "1000110001000111", 15268 => "0101101101001111", 15269 => "0110001010111011", 15270 => "1011001101001111", 15271 => "1011011110110101", 15272 => "1010001000110101", 15273 => "0111001010010010", 15274 => "0110010010111101", 15275 => "1001010110111101", 15276 => "1100001101001011", 15277 => "1110111111101100", 15278 => "1001010000111001", 15279 => "0001000000101101", 15280 => "1101010100101111", 15281 => "1011111001110111", 15282 => "0010110110111101", 15283 => "1010010000100000", 15284 => "0110001110100111", 15285 => "0011110100100010", 15286 => "1110100100010010", 15287 => "1101111101010000", 15288 => "1100010010010111", 15289 => "1101011111000110", 15290 => "0000100000010110", 15291 => "1001001101100001", 15292 => "1001011011000110", 15293 => "0100000101000111", 15294 => "1001001011101100", 15295 => "1110101010011001", 15296 => "1100100011000000", 15297 => "0001110001010100", 15298 => "1010111011000110", 15299 => "1101011001010010", 15300 => "1101010011011110", 15301 => "1000010001101011", 15302 => "0101011110111100", 15303 => "0101010010101101", 15304 => "0100001100100110", 15305 => "0010101110010010", 15306 => "1010011000100010", 15307 => "0100101001011011", 15308 => "0111110110111100", 15309 => "1100110111100000", 15310 => "1000011001111110", 15311 => "1110000101100011", 15312 => "0101001100110011", 15313 => "0000001101011110", 15314 => "1011110111001110", 15315 => "1001011100101010", 15316 => "0011000101010000", 15317 => "1011010000011010", 15318 => "1111110011101110", 15319 => "1000101001111011", 15320 => "1011100110000110", 15321 => "1011011000000010", 15322 => "0101100001111010", 15323 => "1101001011011010", 15324 => "0101110010101100", 15325 => "1111101010101010", 15326 => "0011000000101111", 15327 => "1011101110111111", 15328 => "1010101001001001", 15329 => "0111110111110111", 15330 => "0010100000001011", 15331 => "1110101110001110", 15332 => "1000100011010000", 15333 => "0111100100011001", 15334 => "0111000001100011", 15335 => "0000011000101001", 15336 => "1101111111001010", 15337 => "1000110101000000", 15338 => "1010010001010111", 15339 => "0000010001001011", 15340 => "0010000101001001", 15341 => "1000000101100001", 15342 => "0100011010101100", 15343 => "1111011110010011", 15344 => "0001000111000111", 15345 => "1001110000010000", 15346 => "1010101001101010", 15347 => "1100111000100110", 15348 => "1011011101101111", 15349 => "1111010010001000", 15350 => "0110000001011100", 15351 => "0010011011011001", 15352 => "1010000010001111", 15353 => "1000010000101101", 15354 => "1101011101101101", 15355 => "0000100100100110", 15356 => "1101010101101100", 15357 => "1111000110111011", 15358 => "0111010010110101", 15359 => "1101011111110100", 15360 => "1100111100011101", 15361 => "0011100010000111", 15362 => "0001110101000011", 15363 => "1110111000001011", 15364 => "1010101100110010", 15365 => "0011101100001000", 15366 => "0100000110101101", 15367 => "1101110110001110", 15368 => "1011010000001101", 15369 => "0111011011011010", 15370 => "0101010011011011", 15371 => "1100010111101100", 15372 => "0101111110010111", 15373 => "1100110000111110", 15374 => "1011110101010011", 15375 => "1111010100111100", 15376 => "1001000000101111", 15377 => "0011001100101110", 15378 => "1011011101000110", 15379 => "1001001000000111", 15380 => "0011110011001100", 15381 => "0110001101001001", 15382 => "1101010110101011", 15383 => "1011000111010100", 15384 => "0100111110010101", 15385 => "1001111001101001", 15386 => "1011101001101001", 15387 => "0101010000111110", 15388 => "0100010010111010", 15389 => "0000011011011000", 15390 => "0001000101011100", 15391 => "1001111010001100", 15392 => "1110110111111100", 15393 => "1110011101010110", 15394 => "1100111100001001", 15395 => "1000110100001001", 15396 => "0000000010101101", 15397 => "0000111110101101", 15398 => "0001000000010100", 15399 => "1111001010010110", 15400 => "0110001000100111", 15401 => "0100101111110001", 15402 => "1100010110001010", 15403 => "1000100010101010", 15404 => "1001010001011011", 15405 => "1011100110111010", 15406 => "0000010011110011", 15407 => "1010011001110100", 15408 => "0101011010100111", 15409 => "0110100110111110", 15410 => "0101011110110001", 15411 => "0011110010001111", 15412 => "0000001000110111", 15413 => "1100101011011000", 15414 => "0111100011001011", 15415 => "0010010000011100", 15416 => "1001001111010110", 15417 => "1110001100010011", 15418 => "1100010000000110", 15419 => "0001111001111111", 15420 => "1001010111011000", 15421 => "0011001001111110", 15422 => "1111110000010111", 15423 => "0100011100111010", 15424 => "1110101011010110", 15425 => "1100111001010011", 15426 => "1010100110000010", 15427 => "1011110101101000", 15428 => "0100010010101000", 15429 => "0100111110001111", 15430 => "1100111100101011", 15431 => "0101000000111111", 15432 => "1001000000101010", 15433 => "0100100111011000", 15434 => "0000000101100000", 15435 => "1011000000011001", 15436 => "1001111110000111", 15437 => "1110101010001000", 15438 => "0011100000100011", 15439 => "1101111010000111", 15440 => "0010111011111000", 15441 => "1101111001110110", 15442 => "0010010000100000", 15443 => "1010110011101100", 15444 => "1010100110010111", 15445 => "1101001100100000", 15446 => "1101000000010001", 15447 => "1111000011110001", 15448 => "1011110011101111", 15449 => "0111011001001110", 15450 => "0100111000100111", 15451 => "0010000101011110", 15452 => "1011011011111110", 15453 => "0111010110001011", 15454 => "0000110001111010", 15455 => "0101101101000111", 15456 => "0110010011111011", 15457 => "1000001011010110", 15458 => "1000010101010101", 15459 => "0010111101001000", 15460 => "0101110100011111", 15461 => "1000101000000100", 15462 => "0110000010111100", 15463 => "0111010010011000", 15464 => "0010100000110100", 15465 => "0101001101110001", 15466 => "0100110010000100", 15467 => "1011111001010111", 15468 => "1000101001100111", 15469 => "0011001011100100", 15470 => "1110010100000100", 15471 => "1100011001100100", 15472 => "0101010010011011", 15473 => "1101000110011101", 15474 => "1101100111101111", 15475 => "0010011010010101", 15476 => "1110111110101101", 15477 => "1101011000101110", 15478 => "1001001111010001", 15479 => "0101101000101011", 15480 => "0100111100000011", 15481 => "1011010100100000", 15482 => "1101000110100010", 15483 => "1111110001000111", 15484 => "0111010011000110", 15485 => "1110001110001100", 15486 => "0010010001010111", 15487 => "0011011101011111", 15488 => "1011011000100011", 15489 => "0101100001101101", 15490 => "1110001111110101", 15491 => "0001001101100001", 15492 => "1100001100010101", 15493 => "1101000000111111", 15494 => "0110110011111011", 15495 => "0101100000010000", 15496 => "0101101000010111", 15497 => "1010110111011100", 15498 => "0011110110101111", 15499 => "0101011010010110", 15500 => "0101100110011110", 15501 => "1000001111011101", 15502 => "0110010000111111", 15503 => "0011100001111001", 15504 => "1011000011100011", 15505 => "1101100111100001", 15506 => "1100110011110101", 15507 => "0100110111001000", 15508 => "1110001101100100", 15509 => "0111000110110011", 15510 => "0001011010011100", 15511 => "0010000011010101", 15512 => "1011011110110011", 15513 => "0111110101010010", 15514 => "1111110001000010", 15515 => "0000110100001101", 15516 => "1001101101010100", 15517 => "1111010001101101", 15518 => "0001010011101000", 15519 => "0101010001011100", 15520 => "0100110001101101", 15521 => "0010111001100010", 15522 => "0011011100000100", 15523 => "0000010100000100", 15524 => "0001000001110100", 15525 => "0100101100110010", 15526 => "1001111010101000", 15527 => "1011101101011101", 15528 => "1000101010010100", 15529 => "1101100111100001", 15530 => "1111111110011110", 15531 => "1011111111001110", 15532 => "1110101010110111", 15533 => "1110100010001000", 15534 => "0110110011101110", 15535 => "0001001010101100", 15536 => "0100000100011010", 15537 => "1000001110101001", 15538 => "1111110111110111", 15539 => "1110101000111000", 15540 => "0010111100100110", 15541 => "0110001111011010", 15542 => "0001111000111100", 15543 => "1101011001000001", 15544 => "1011111110001001", 15545 => "1011011101001101", 15546 => "1000101001101001", 15547 => "1011100011000100", 15548 => "0100101001100101", 15549 => "1100100111100000", 15550 => "0100100011111111", 15551 => "0100010010001011", 15552 => "1100011011001100", 15553 => "0110111111111100", 15554 => "1000101010010000", 15555 => "1010100000010101", 15556 => "1011110101001000", 15557 => "0111111010111001", 15558 => "0010111011011101", 15559 => "1101110100001101", 15560 => "1010111000010010", 15561 => "0101011001100011", 15562 => "0001101001000001", 15563 => "0100011010101100", 15564 => "1101010010111011", 15565 => "1100100000110110", 15566 => "0101111110000011", 15567 => "1011011101000010", 15568 => "0000011001000001", 15569 => "0000000001001101", 15570 => "1100110010110110", 15571 => "1010110000111011", 15572 => "0101101111010100", 15573 => "1101001101100100", 15574 => "0001001011001101", 15575 => "0101101100101110", 15576 => "0001010101001001", 15577 => "0110011000011000", 15578 => "0111001000000000", 15579 => "1001000010111111", 15580 => "1001110011100011", 15581 => "1000100101110001", 15582 => "1111110011100111", 15583 => "1011001100011001", 15584 => "1110010101110101", 15585 => "0011000000010011", 15586 => "0110100111101011", 15587 => "0101100010000001", 15588 => "1010000111100101", 15589 => "0000111110000111", 15590 => "1111011100100001", 15591 => "0011000011010111", 15592 => "0001100010011000", 15593 => "1110011100010011", 15594 => "0111011000101111", 15595 => "1011110010110010", 15596 => "0010110010110101", 15597 => "1101110100011101", 15598 => "1111111111010101", 15599 => "0110111110000011", 15600 => "1010001010011111", 15601 => "1111010010001011", 15602 => "1010011100011100", 15603 => "1010001111011101", 15604 => "0000011000010101", 15605 => "1111011110011101", 15606 => "0110001011000111", 15607 => "0100101001111010", 15608 => "0100011011110100", 15609 => "0100011011001111", 15610 => "1000011001101110", 15611 => "1100001000011111", 15612 => "0011001010010101", 15613 => "0101010000100010", 15614 => "0100001101110010", 15615 => "1011000001111101", 15616 => "1111111100011010", 15617 => "1100011111001101", 15618 => "0100000101110011", 15619 => "1001101000111111", 15620 => "0001001010100111", 15621 => "1000000010001011", 15622 => "1110010111110101", 15623 => "0111011100111001", 15624 => "0011101011111000", 15625 => "0011110101100000", 15626 => "0001000100000110", 15627 => "0110001000100000", 15628 => "0100010011000001", 15629 => "1001100100100010", 15630 => "1110101001100001", 15631 => "1110111010001100", 15632 => "0101011010001100", 15633 => "1110101010111100", 15634 => "1100001001001011", 15635 => "0101110011000101", 15636 => "1010100100011001", 15637 => "1101111011001100", 15638 => "1010100011100010", 15639 => "1111001100101100", 15640 => "0011011010111010", 15641 => "0101111000101101", 15642 => "0111001111001000", 15643 => "1001010100100101", 15644 => "0011100101001110", 15645 => "1000001011011111", 15646 => "1110101000010111", 15647 => "0001100001111100", 15648 => "0000010111000100", 15649 => "0101110001000101", 15650 => "0101011000000111", 15651 => "1001010001100000", 15652 => "0010000000000101", 15653 => "0111110010100001", 15654 => "1101100111111100", 15655 => "1010001011110100", 15656 => "1001111100010111", 15657 => "0010010101101100", 15658 => "0101001110000011", 15659 => "1110011110000110", 15660 => "1000001000001011", 15661 => "0111000000100111", 15662 => "0010101110110000", 15663 => "0101111111001101", 15664 => "1111101000101101", 15665 => "1111000011110110", 15666 => "0100111100111101", 15667 => "0110011000000100", 15668 => "0101001001111011", 15669 => "1100010110110010", 15670 => "0111110011101000", 15671 => "1101001111001001", 15672 => "0110110110001110", 15673 => "0010111011110110", 15674 => "1011111101010010", 15675 => "1110001111101011", 15676 => "0011000110110000", 15677 => "0100101010111011", 15678 => "0000111010100001", 15679 => "1000111001111001", 15680 => "0101011111111000", 15681 => "1010111101101110", 15682 => "1101010111111011", 15683 => "0001001100101100", 15684 => "1011110111011011", 15685 => "0111111111101101", 15686 => "1010010001001110", 15687 => "0100111101100110", 15688 => "1001000011011111", 15689 => "0100111110010111", 15690 => "1011110101010010", 15691 => "0001011010111111", 15692 => "0101000010100011", 15693 => "0001101000000001", 15694 => "0010110011100011", 15695 => "1110101011000100", 15696 => "1010101111011100", 15697 => "0001001001100000", 15698 => "1101111100101111", 15699 => "0101000000100011", 15700 => "0010111101100010", 15701 => "0000101101111111", 15702 => "1001011100010011", 15703 => "0100000001110010", 15704 => "0010101111001111", 15705 => "0111110101111010", 15706 => "1011000000100111", 15707 => "1111010000101101", 15708 => "0101011001110001", 15709 => "1101110010000111", 15710 => "0111100001111111", 15711 => "1101110001011101", 15712 => "1100110000000011", 15713 => "1100111001110100", 15714 => "0010010110001000", 15715 => "1111000010010110", 15716 => "0110001101010111", 15717 => "1011100001111011", 15718 => "0111011011111000", 15719 => "1110001101010000", 15720 => "1101101100001011", 15721 => "1111011110001101", 15722 => "0101010100000001", 15723 => "1010010001110000", 15724 => "0111100010010110", 15725 => "1000100100001111", 15726 => "0101101011101111", 15727 => "1011011110101011", 15728 => "1011100011000010", 15729 => "0110111001110001", 15730 => "0001000110111011", 15731 => "1000010001101101", 15732 => "1100101100111010", 15733 => "0000010001000011", 15734 => "1011100110111011", 15735 => "1000110111000101", 15736 => "0101101110000101", 15737 => "0011100110000111", 15738 => "0011110110100110", 15739 => "1110110010011010", 15740 => "1101110011010011", 15741 => "1010001101010011", 15742 => "0000000001100111", 15743 => "1100111011000000", 15744 => "1101001100010001", 15745 => "0011011101001010", 15746 => "1110000111110101", 15747 => "0101110001011101", 15748 => "1000110101101011", 15749 => "1110110001111100", 15750 => "1001000110100001", 15751 => "1001001100000011", 15752 => "0100110111110000", 15753 => "0000001011111011", 15754 => "1101001011111010", 15755 => "0101011000011011", 15756 => "0111111001101111", 15757 => "1110010100111001", 15758 => "0001111110111111", 15759 => "0000100110011000", 15760 => "1010110100100111", 15761 => "1111101001100010", 15762 => "1111100000100000", 15763 => "1000101000000111", 15764 => "1110011110011010", 15765 => "0011110000001010", 15766 => "0100111101110111", 15767 => "1011011101110010", 15768 => "0011000101101111", 15769 => "1011110101110010", 15770 => "0101100101000010", 15771 => "0011000100111100", 15772 => "1011000110000100", 15773 => "1010111101100111", 15774 => "1010110100101110", 15775 => "0100011001111000", 15776 => "1000111010011110", 15777 => "1011000100100111", 15778 => "1011111000111001", 15779 => "1101111001001110", 15780 => "1101100000011100", 15781 => "1100011101010010", 15782 => "1010110000110111", 15783 => "0000011000011100", 15784 => "1110100011100011", 15785 => "1000111000110101", 15786 => "0100111000011110", 15787 => "0100010010000111", 15788 => "0110010110010101", 15789 => "1000111011010010", 15790 => "1000011111000100", 15791 => "0110010111110000", 15792 => "0111000110100010", 15793 => "0110100011010000", 15794 => "0110000100110011", 15795 => "0010111101011110", 15796 => "1001110101110101", 15797 => "0101010000000101", 15798 => "1010100111111110", 15799 => "1001001010011000", 15800 => "0101011000100100", 15801 => "0010111001100001", 15802 => "0001100001001111", 15803 => "1011111101101111", 15804 => "0110111100101001", 15805 => "1111101111010011", 15806 => "1000011111110101", 15807 => "0000010111000001", 15808 => "0011110000011100", 15809 => "0110101010111011", 15810 => "1010100101001100", 15811 => "1110000000110111", 15812 => "0000011001001101", 15813 => "1011000000101010", 15814 => "1010111010000101", 15815 => "0110101110011100", 15816 => "0100101101111110", 15817 => "0101101010101010", 15818 => "0110011010001100", 15819 => "0111001101111000", 15820 => "0111001100010110", 15821 => "1110110001110000", 15822 => "0001110111111110", 15823 => "0010111010010001", 15824 => "0101110011011001", 15825 => "0111011100100011", 15826 => "1110101000101111", 15827 => "0000101001001011", 15828 => "0110001100110000", 15829 => "0111101010011101", 15830 => "1111000100010100", 15831 => "1100111101100001", 15832 => "0100101111111010", 15833 => "1010010011110000", 15834 => "0001001011001111", 15835 => "1100110110101110", 15836 => "1110111010011000", 15837 => "0110010101011100", 15838 => "0011010011101001", 15839 => "1101111011011111", 15840 => "1101001011001000", 15841 => "1000111010011110", 15842 => "0100100001001000", 15843 => "0001100101100100", 15844 => "0011110000110100", 15845 => "0000001110010011", 15846 => "0101000000001110", 15847 => "0110111011101100", 15848 => "1010000011101000", 15849 => "1011101000110100", 15850 => "1011110100001100", 15851 => "1001111010101101", 15852 => "1111100010101110", 15853 => "1000001100101001", 15854 => "1000100011001110", 15855 => "1101101001011101", 15856 => "0000110101010110", 15857 => "0000110011110010", 15858 => "1110010010101000", 15859 => "0111110011000101", 15860 => "0011110111000110", 15861 => "0101110100101011", 15862 => "0100100001101000", 15863 => "0001101011001100", 15864 => "0010011000001001", 15865 => "1100111010011110", 15866 => "1011001011011000", 15867 => "0110001010110100", 15868 => "1101101010111001", 15869 => "0111001101101011", 15870 => "0001110101011100", 15871 => "1111001100011110", 15872 => "1010110010110001", 15873 => "1100011101101100", 15874 => "1110111000011100", 15875 => "0111110110111010", 15876 => "1111000000010010", 15877 => "1010111011110011", 15878 => "0110000011111001", 15879 => "1111100001001010", 15880 => "0000110101101000", 15881 => "0100100100010001", 15882 => "1101111010110011", 15883 => "0100101111000001", 15884 => "0101100101110011", 15885 => "1001000101001001", 15886 => "0100101111111111", 15887 => "1011110101101010", 15888 => "1001100101100111", 15889 => "1110011100011110", 15890 => "1100010110110001", 15891 => "1000011100001110", 15892 => "1011100000100001", 15893 => "0110010101100000", 15894 => "1111001111101111", 15895 => "1000111000111111", 15896 => "0010110011001111", 15897 => "0111011001101110", 15898 => "0011100011111011", 15899 => "0111001011011000", 15900 => "0100000011100110", 15901 => "0010000000011001", 15902 => "1001000000110000", 15903 => "1000010101110001", 15904 => "1101000001011010", 15905 => "1010000000010000", 15906 => "0101101110100101", 15907 => "0000011110000010", 15908 => "1001011101101101", 15909 => "1110011111011100", 15910 => "1011000001010111", 15911 => "0111011111100010", 15912 => "1001011011000000", 15913 => "0111100101110100", 15914 => "1001111101000111", 15915 => "1010010100101111", 15916 => "1100011010001111", 15917 => "1100011110100011", 15918 => "0110110010110000", 15919 => "0000010000101111", 15920 => "1000001000000000", 15921 => "0000010101100111", 15922 => "1010100011001100", 15923 => "1100111100001001", 15924 => "1100111101011111", 15925 => "1111011101100110", 15926 => "0111100011111001", 15927 => "0101110110011000", 15928 => "0000001101110101", 15929 => "0001111110010001", 15930 => "1000011100010100", 15931 => "1111100100110100", 15932 => "1000010110011110", 15933 => "0100001101011001", 15934 => "1101001111000111", 15935 => "1101101101010110", 15936 => "1011101010101010", 15937 => "1001001000101001", 15938 => "0101001000001010", 15939 => "0010010111000001", 15940 => "0101101011111110", 15941 => "1001110001111001", 15942 => "1001001000111111", 15943 => "1000111011001001", 15944 => "0000100111100111", 15945 => "1110101000011011", 15946 => "1010100101110110", 15947 => "0110100110011101", 15948 => "1010011110111111", 15949 => "0100111111110011", 15950 => "0101011111101011", 15951 => "1001001110000001", 15952 => "0110110011001001", 15953 => "1101111000000111", 15954 => "1110111000010001", 15955 => "0011100100111011", 15956 => "0101111100100001", 15957 => "1001001100001101", 15958 => "0100110101010011", 15959 => "1011100000010001", 15960 => "0101100100111100", 15961 => "0101011101010011", 15962 => "0001110001001010", 15963 => "0011110000011010", 15964 => "1010111011111010", 15965 => "0111101110101000", 15966 => "0000000111010011", 15967 => "0110101011011010", 15968 => "1010011101011011", 15969 => "0010010001000111", 15970 => "1011110000101100", 15971 => "0101111010111011", 15972 => "0001111011011101", 15973 => "1101000101000001", 15974 => "0000000111101010", 15975 => "0010111000010000", 15976 => "1011110110101001", 15977 => "0101000000001110", 15978 => "0011011001010110", 15979 => "1101110111101011", 15980 => "0100000010011101", 15981 => "0011100111001110", 15982 => "0101101000000001", 15983 => "1101001101010110", 15984 => "0000101010110111", 15985 => "0011110111110011", 15986 => "1001100110110101", 15987 => "0010000010110111", 15988 => "1010111000111001", 15989 => "0000000001001000", 15990 => "0011011010111100", 15991 => "1000001010011000", 15992 => "1000001001100101", 15993 => "1100100011000100", 15994 => "1001111100000100", 15995 => "1111011000100000", 15996 => "0101001010111111", 15997 => "1110111111100011", 15998 => "0111011000001110", 15999 => "0101101101001000", 16000 => "1101110101110010", 16001 => "1010011111001100", 16002 => "0100100011000001", 16003 => "0000110100000010", 16004 => "1001100110111000", 16005 => "1010010011110010", 16006 => "0101101110001001", 16007 => "0010001000010011", 16008 => "1111101011100110", 16009 => "0000111000100011", 16010 => "1011110100011100", 16011 => "0100101011110111", 16012 => "1110101111110100", 16013 => "0010010111001110", 16014 => "1001110111100001", 16015 => "1000101001110100", 16016 => "0010111000101010", 16017 => "0000111000011001", 16018 => "0100010111010101", 16019 => "1011110010101011", 16020 => "0111100101111001", 16021 => "1011101100001011", 16022 => "0110001111100001", 16023 => "0011101101011011", 16024 => "0111110100100001", 16025 => "1110010110000001", 16026 => "0010111011000100", 16027 => "0000100100001010", 16028 => "1111000110101101", 16029 => "1111011101110100", 16030 => "0000110011000001", 16031 => "1100001100110100", 16032 => "1110111101010010", 16033 => "0011000000110010", 16034 => "1000010001001011", 16035 => "0010110000010011", 16036 => "1000001101010011", 16037 => "1100101111110011", 16038 => "1110100010011111", 16039 => "1110000010000100", 16040 => "1011100100110111", 16041 => "1001000110100101", 16042 => "0101111011101110", 16043 => "1111010000011111", 16044 => "1010100001000011", 16045 => "0001100101000110", 16046 => "0000100010110111", 16047 => "0100101101010011", 16048 => "1001111000011100", 16049 => "1101010100000000", 16050 => "1111000111111011", 16051 => "1100100010110001", 16052 => "1111000011011010", 16053 => "1011101110100010", 16054 => "0110010111110000", 16055 => "1010111011100110", 16056 => "1111000101111100", 16057 => "0011001010111010", 16058 => "0010001101010000", 16059 => "1100000100110011", 16060 => "0001000110110011", 16061 => "1000111000000011", 16062 => "1111000010000100", 16063 => "1011000011001111", 16064 => "1101001110101011", 16065 => "0000000010110001", 16066 => "0110011100001001", 16067 => "0001001111100101", 16068 => "0011011100111111", 16069 => "1100110010111100", 16070 => "1010000011011010", 16071 => "1110110111111010", 16072 => "0111000111001111", 16073 => "1011111001000011", 16074 => "1001101011100100", 16075 => "0010010111100010", 16076 => "0010100000101100", 16077 => "0111001000011110", 16078 => "0101111100101100", 16079 => "0111010000100101", 16080 => "0100111111011101", 16081 => "1111010010101010", 16082 => "0111100010000100", 16083 => "0010010010101101", 16084 => "1010001010110011", 16085 => "0101001111111010", 16086 => "1100010010010011", 16087 => "0000011110011010", 16088 => "0100011111000100", 16089 => "0000101100000010", 16090 => "1001001001101000", 16091 => "0101001101010010", 16092 => "0100010010000110", 16093 => "1100000011100010", 16094 => "1011000010011000", 16095 => "1010111010000111", 16096 => "1001100111100000", 16097 => "0010010010010100", 16098 => "1110010110010111", 16099 => "0101010111111111", 16100 => "0111110110101111", 16101 => "1010110111001011", 16102 => "1000100000001001", 16103 => "1000011100001010", 16104 => "1011110011111100", 16105 => "1100111000011101", 16106 => "1111100111111001", 16107 => "1110100110011010", 16108 => "1110100110110100", 16109 => "0110000001100101", 16110 => "1001000001100111", 16111 => "1011001100001110", 16112 => "0001001010111110", 16113 => "0001010000110001", 16114 => "1101011101100100", 16115 => "1011110101111011", 16116 => "1100110000110101", 16117 => "0010000000010111", 16118 => "1100110000011000", 16119 => "1110101001000001", 16120 => "0001111100111111", 16121 => "1010111000101100", 16122 => "1110011001100100", 16123 => "0110011111010001", 16124 => "1111011111111001", 16125 => "0011111000011111", 16126 => "1010111011111111", 16127 => "1110110001001010", 16128 => "1110000111110010", 16129 => "1111100011101111", 16130 => "1110101011011110", 16131 => "0001010010010011", 16132 => "0001010001110001", 16133 => "0011100000110110", 16134 => "1111101000000100", 16135 => "0110100010010111", 16136 => "0101001000111110", 16137 => "0010110011000110", 16138 => "0110111110110100", 16139 => "0110001011111010", 16140 => "1011011100101001", 16141 => "0001101111100011", 16142 => "0001100001111110", 16143 => "1110111101000011", 16144 => "0111011101100001", 16145 => "1100110101000010", 16146 => "1010011110010101", 16147 => "1001100100101101", 16148 => "0000001111010111", 16149 => "1011110100011000", 16150 => "0100111010010010", 16151 => "1000101101100001", 16152 => "1000110000001111", 16153 => "0011000011110001", 16154 => "0010110010100010", 16155 => "0000000010100101", 16156 => "1111111111001110", 16157 => "1111010010000101", 16158 => "1010110011101111", 16159 => "0100010100101001", 16160 => "0011001010111011", 16161 => "1011101100000110", 16162 => "1001011001010010", 16163 => "0111110000001011", 16164 => "1110100110111111", 16165 => "1010101110101010", 16166 => "0010010110111111", 16167 => "0100010110100011", 16168 => "1000000001011011", 16169 => "1100111010011100", 16170 => "0000011001010110", 16171 => "1011011101100100", 16172 => "1111111101100111", 16173 => "1101000000001011", 16174 => "0100010110101111", 16175 => "0111001100101000", 16176 => "0111001110010000", 16177 => "1110110000110101", 16178 => "1001001100000001", 16179 => "1010011011011101", 16180 => "0111011101010001", 16181 => "1010100101001110", 16182 => "1000010110111101", 16183 => "0000010110111111", 16184 => "0101110011101101", 16185 => "0101001110100110", 16186 => "1000001001011011", 16187 => "1001111001111001", 16188 => "0110110101111101", 16189 => "0000000000011110", 16190 => "1110011111001111", 16191 => "1100011111000011", 16192 => "1100101100011001", 16193 => "0111101010111111", 16194 => "0000011001100101", 16195 => "1110100110111100", 16196 => "0101111011100001", 16197 => "0011100001111100", 16198 => "0001101000111001", 16199 => "0001000011010111", 16200 => "1000010110101101", 16201 => "1011101011011010", 16202 => "0001100001001100", 16203 => "1111011010100111", 16204 => "1010100111111110", 16205 => "1011111100000101", 16206 => "0001010100000111", 16207 => "1111101000101011", 16208 => "1101110111100110", 16209 => "1011011110001101", 16210 => "0011000001001010", 16211 => "0110010000110111", 16212 => "0001000001111110", 16213 => "0101100000111100", 16214 => "0100001011101110", 16215 => "1101011101100001", 16216 => "0000101110110101", 16217 => "1000000011010111", 16218 => "1000111011101001", 16219 => "0101110000100110", 16220 => "0010100010111100", 16221 => "1110000000000111", 16222 => "1101010101010101", 16223 => "1110000110001011", 16224 => "1101000110000100", 16225 => "1110100101100010", 16226 => "0011101111010110", 16227 => "0111101000011001", 16228 => "1011000000101000", 16229 => "1010101111011110", 16230 => "1001001010000011", 16231 => "1000100001001100", 16232 => "0010000000010101", 16233 => "0101111010011111", 16234 => "0100011011111011", 16235 => "1100011100111100", 16236 => "0000100111100000", 16237 => "0010100011110111", 16238 => "1000100010110000", 16239 => "1010100011110010", 16240 => "1001100001000100", 16241 => "1100101100000010", 16242 => "0011110110111101", 16243 => "1100000111000011", 16244 => "0011000011010110", 16245 => "1100010110100000", 16246 => "0001110000110111", 16247 => "1111000011000101", 16248 => "1010101010000100", 16249 => "1110011101000111", 16250 => "1111101100001101", 16251 => "0111110011100010", 16252 => "1110110100101001", 16253 => "1010101001100011", 16254 => "0001101010010111", 16255 => "0111010001110111", 16256 => "1000100101110100", 16257 => "1011010111010001", 16258 => "1000000011010100", 16259 => "1101001100011011", 16260 => "0001111111101011", 16261 => "1000100110101110", 16262 => "0010000000101000", 16263 => "1100111000011010", 16264 => "0000010010001110", 16265 => "0001100101111100", 16266 => "1010011110000110", 16267 => "1000000000010111", 16268 => "1110011101001011", 16269 => "1111111110110110", 16270 => "0000000111010010", 16271 => "0010000000001001", 16272 => "0100011101010110", 16273 => "0010100001001111", 16274 => "1111010001111010", 16275 => "0000000011110000", 16276 => "1110100000011010", 16277 => "0011110001101110", 16278 => "1110000010010110", 16279 => "0100001010111110", 16280 => "1000101101011100", 16281 => "1110010001011110", 16282 => "1010111001110101", 16283 => "1111001010000011", 16284 => "0010100000010110", 16285 => "0111101001011001", 16286 => "0100011001001100", 16287 => "0000111101110110", 16288 => "0011010011101101", 16289 => "0001101001110110", 16290 => "1011110000110001", 16291 => "1001010101100110", 16292 => "0111011010011011", 16293 => "1101101110011101", 16294 => "1111011110110001", 16295 => "1001110100011011", 16296 => "0010010000010011", 16297 => "0011000100001101", 16298 => "0011001100010110", 16299 => "1110101011000011", 16300 => "1011011000110110", 16301 => "0000111101101100", 16302 => "0011100000101100", 16303 => "0100101010111110", 16304 => "0000010100011011", 16305 => "1000101101010100", 16306 => "0100010011000110", 16307 => "0001000110011001", 16308 => "1110011110011100", 16309 => "1110110000110011", 16310 => "1001001001101011", 16311 => "0111111000100111", 16312 => "1110000101011000", 16313 => "1010111111010110", 16314 => "1110100110101101", 16315 => "1010101111101011", 16316 => "0000011110110011", 16317 => "1000000011100111", 16318 => "0110000101101111", 16319 => "1000000110110010", 16320 => "1111110100001010", 16321 => "1111100100111110", 16322 => "0100101111001101", 16323 => "0001011001100010", 16324 => "0010011101001110", 16325 => "0001111111101100", 16326 => "0101000011100011", 16327 => "1001111101101100", 16328 => "0010101000101011", 16329 => "1100110001110110", 16330 => "0011100000001001", 16331 => "1001100110110001", 16332 => "1001111010001111", 16333 => "1100100101001110", 16334 => "1000110010001010", 16335 => "0011111001100000", 16336 => "1101100110100000", 16337 => "0110101011110110", 16338 => "0111111010110101", 16339 => "1000101000101001", 16340 => "0000000001010001", 16341 => "0001100011111100", 16342 => "1100000100100101", 16343 => "1011001111011110", 16344 => "1100001010100100", 16345 => "0100010100011011", 16346 => "1101000111110110", 16347 => "1011101001100010", 16348 => "0010110011010100", 16349 => "0111001111010110", 16350 => "0010110001110011", 16351 => "1111100001110011", 16352 => "0001100000000110", 16353 => "0010011000111110", 16354 => "0000111100001111", 16355 => "0000000101010111", 16356 => "1111101100101001", 16357 => "1000001010100100", 16358 => "0111101011101100", 16359 => "1101101100100010", 16360 => "0101011100100100", 16361 => "1111001101000101", 16362 => "1100010000011001", 16363 => "1010100011101101", 16364 => "1001101111110001", 16365 => "1001110011100101", 16366 => "1110101001101001", 16367 => "0000111011111110", 16368 => "1110111101011100", 16369 => "0011010101001000", 16370 => "1100001100010111", 16371 => "1001011001111110", 16372 => "1011000010101101", 16373 => "1101000111000101", 16374 => "1111001101001000", 16375 => "1110110110110001", 16376 => "0011101110110001", 16377 => "0100011101000011", 16378 => "1111101010011011", 16379 => "0101111101001110", 16380 => "0111000100011001", 16381 => "0000000011100000", 16382 => "1101000010100000", 16383 => "0000100000000000", 16384 => "1010101101110101", 16385 => "1010101001001110", 16386 => "0110100011110110", 16387 => "0010001010000001", 16388 => "1001000011011111", 16389 => "0111110011110001", 16390 => "1110010111110010", 16391 => "1101001000100010", 16392 => "1110000100000010", 16393 => "1101100111010111", 16394 => "1011011000010111", 16395 => "1000101101000000", 16396 => "0010110100100110", 16397 => "0001101111111111", 16398 => "1000111110000110", 16399 => "0010111111001111", 16400 => "1001001010110101", 16401 => "0011110111100101", 16402 => "0010101000000110", 16403 => "1000001001011001", 16404 => "0110000100110110", 16405 => "0110111100000100", 16406 => "1011000100100100", 16407 => "1011101110001100", 16408 => "0110111110001111", 16409 => "1110100010110100", 16410 => "0101101011111101", 16411 => "1001101011100001", 16412 => "0000000110001010", 16413 => "1000011110110111", 16414 => "0001101111010101", 16415 => "0001011111001110", 16416 => "1100010010101000", 16417 => "0010000101001110", 16418 => "0011100011000001", 16419 => "1010100010010111", 16420 => "1000001110111101", 16421 => "0100100101011101", 16422 => "0001001110000110", 16423 => "0111111010000000", 16424 => "1111101011000101", 16425 => "1110101000110101", 16426 => "0001001001110001", 16427 => "0111010011000010", 16428 => "0110001111110000", 16429 => "1011110000000110", 16430 => "0000101101111001", 16431 => "0001010100111011", 16432 => "1010010101010101", 16433 => "1100110010000111", 16434 => "0110000101111010", 16435 => "1011000101011010", 16436 => "1000000101101101", 16437 => "0000101000100100", 16438 => "1001111100010100", 16439 => "0010110110101001", 16440 => "0110000111110011", 16441 => "0010110000111100", 16442 => "0000110001001111", 16443 => "0011001000101101", 16444 => "0010011101011011", 16445 => "0101010010101111", 16446 => "0011010010001101", 16447 => "1111110100111001", 16448 => "0100111100101011", 16449 => "0111010010101111", 16450 => "0111100011011101", 16451 => "0001000000111010", 16452 => "0101010000001011", 16453 => "1001001110100000", 16454 => "1100101101111111", 16455 => "1010100011011101", 16456 => "1111101000110111", 16457 => "0110000010011110", 16458 => "0110111000011100", 16459 => "1000101001000111", 16460 => "0101101100000010", 16461 => "0111011000010001", 16462 => "0111010111101011", 16463 => "1000000001000100", 16464 => "1010011011011111", 16465 => "0011011010000111", 16466 => "1010011110010000", 16467 => "1110111011001011", 16468 => "0011000100100110", 16469 => "1111111010001101", 16470 => "0010101010110001", 16471 => "1001001010000101", 16472 => "1101011101111001", 16473 => "0100010110000001", 16474 => "0100011100000110", 16475 => "1010001100101011", 16476 => "0010111100101100", 16477 => "0111110000111111", 16478 => "1110101011110100", 16479 => "1100100110011111", 16480 => "0111001010010011", 16481 => "0111111010101101", 16482 => "0110010001100110", 16483 => "1110011100001000", 16484 => "1000001111000001", 16485 => "1101111101010110", 16486 => "0010011110110101", 16487 => "0100010110100011", 16488 => "0011011000011011", 16489 => "1100011110011010", 16490 => "1001111010000010", 16491 => "0111001011011010", 16492 => "0011100001101111", 16493 => "0010100000100001", 16494 => "0110001010011111", 16495 => "1001010000111000", 16496 => "1111001010110110", 16497 => "0011110000101000", 16498 => "1110000000001001", 16499 => "1100111101000001", 16500 => "1010010011110000", 16501 => "0011100111001110", 16502 => "0011011010001111", 16503 => "1011010111000011", 16504 => "1011111101011110", 16505 => "0100010100001001", 16506 => "1011011100100001", 16507 => "0110111011001101", 16508 => "1000110110101010", 16509 => "1100100011111111", 16510 => "0110011101110111", 16511 => "0101111000101001", 16512 => "1010111011010111", 16513 => "1111111111100101", 16514 => "0010100101101001", 16515 => "0110111011100000", 16516 => "1111111111000110", 16517 => "0111001000000000", 16518 => "0001000101111000", 16519 => "1110010100000110", 16520 => "0010110000011110", 16521 => "0001011011110100", 16522 => "1010001001001111", 16523 => "0110001111110101", 16524 => "0111100110100101", 16525 => "1010011101100001", 16526 => "1001101001110111", 16527 => "0010011110001011", 16528 => "0000110111110100", 16529 => "0001100011110111", 16530 => "1010011100100110", 16531 => "1110011100111101", 16532 => "0100001010010101", 16533 => "0000011010100000", 16534 => "0011011100111010", 16535 => "1101010111001011", 16536 => "0001010111101110", 16537 => "1011101111000001", 16538 => "1010010011010000", 16539 => "0110001001001110", 16540 => "1000001010101000", 16541 => "1110110001110111", 16542 => "1000010000000000", 16543 => "1111100000010011", 16544 => "0001001001100001", 16545 => "0001100001100000", 16546 => "0100110101111001", 16547 => "0111100111000110", 16548 => "1001010001000011", 16549 => "1111110110110010", 16550 => "0111111000001100", 16551 => "1010101111110010", 16552 => "0100101001001100", 16553 => "0001101010100000", 16554 => "0101001100111100", 16555 => "0000101011101101", 16556 => "0101010001001110", 16557 => "0100101101100101", 16558 => "0110111010011110", 16559 => "1011110010001100", 16560 => "0111000101000000", 16561 => "0101111110001101", 16562 => "0100111111100010", 16563 => "0101001000000110", 16564 => "1110010111111001", 16565 => "1111011101100111", 16566 => "0001100101010111", 16567 => "1000111101011000", 16568 => "1011011100011001", 16569 => "0100000011011000", 16570 => "0110000011100110", 16571 => "0001111011110000", 16572 => "0001101110000100", 16573 => "1011111011010101", 16574 => "0111101010110111", 16575 => "1111100011001000", 16576 => "1011000111000001", 16577 => "1101100010000000", 16578 => "1001100011100110", 16579 => "0010111011011110", 16580 => "0110100110110011", 16581 => "1010011101111001", 16582 => "1111011000011010", 16583 => "0101011111111100", 16584 => "1011010101111010", 16585 => "0110000001001101", 16586 => "0010000111101010", 16587 => "0010000000101010", 16588 => "1011000010001010", 16589 => "1111110001011110", 16590 => "0110000100111011", 16591 => "0100000001101011", 16592 => "0001101000000101", 16593 => "0000000000001110", 16594 => "1000111010001010", 16595 => "1000111100001000", 16596 => "1111101001101010", 16597 => "0110001001100000", 16598 => "1000111011001101", 16599 => "0111111110110010", 16600 => "0000000010101100", 16601 => "1110001111000010", 16602 => "1100000111000101", 16603 => "1010111000000000", 16604 => "0111111100000010", 16605 => "0100110010001010", 16606 => "0101000000111001", 16607 => "1010111101000010", 16608 => "1100111101110101", 16609 => "0010110101001000", 16610 => "0000100111100000", 16611 => "0011000010110000", 16612 => "0110011001001011", 16613 => "0010111011100001", 16614 => "1110111000100010", 16615 => "1111000110100100", 16616 => "1101010011001011", 16617 => "0111101001010000", 16618 => "0010100101000011", 16619 => "1101101011100001", 16620 => "1010111011110011", 16621 => "0101100001010001", 16622 => "1011111100110000", 16623 => "1000100110010001", 16624 => "1101000001000101", 16625 => "0000101001010000", 16626 => "0111000101100000", 16627 => "1111000001000110", 16628 => "1101011110100001", 16629 => "1110001010100111", 16630 => "0101100011001111", 16631 => "1101010111111000", 16632 => "0101110000001100", 16633 => "0110010110101000", 16634 => "1101110011001010", 16635 => "1101001011010111", 16636 => "1100001000011101", 16637 => "0111101101011110", 16638 => "1000101011011010", 16639 => "1010010110100110", 16640 => "0100101001111101", 16641 => "0001100010101101", 16642 => "1001011001111110", 16643 => "0010000001000001", 16644 => "0001000011011100", 16645 => "1001101000100101", 16646 => "1000000010011100", 16647 => "1101101011100000", 16648 => "1000000001101010", 16649 => "0000111001110101", 16650 => "1101100101100011", 16651 => "0010011010110110", 16652 => "1011000010100011", 16653 => "0000001101010011", 16654 => "1100000110100011", 16655 => "0100010101011011", 16656 => "0110011011111111", 16657 => "1110100011101010", 16658 => "0000011100010000", 16659 => "0100010101111010", 16660 => "1010001011001010", 16661 => "1011010111111001", 16662 => "0000011011100000", 16663 => "0001111110111010", 16664 => "1010101111111101", 16665 => "0110110101111000", 16666 => "1111011111000001", 16667 => "1110011010100011", 16668 => "0110100111110001", 16669 => "0101010100010010", 16670 => "1000111110001011", 16671 => "1110110010110111", 16672 => "0101101011010111", 16673 => "0110110111000100", 16674 => "0000011011010001", 16675 => "0010100010110011", 16676 => "0101001101010000", 16677 => "1001111100100001", 16678 => "1010100000111000", 16679 => "1011110011110011", 16680 => "0000010110111000", 16681 => "1100101101110111", 16682 => "0000010111011011", 16683 => "0101010001001111", 16684 => "1001111010101010", 16685 => "1101101111000101", 16686 => "1001101011101000", 16687 => "0010010001011001", 16688 => "0010010110100011", 16689 => "1011000111010001", 16690 => "1011010100110010", 16691 => "1000111010100010", 16692 => "1011000111100100", 16693 => "1101010011010100", 16694 => "1011100101011011", 16695 => "0001101000011011", 16696 => "1101000110010100", 16697 => "1100110011111010", 16698 => "1101101000110101", 16699 => "0010001110011110", 16700 => "1101100110000011", 16701 => "1000111011001100", 16702 => "1010010110100101", 16703 => "1000000000000000", 16704 => "0000101100110111", 16705 => "1101010011110101", 16706 => "1000010110100000", 16707 => "1110111010111100", 16708 => "0010001111100101", 16709 => "1111100010011100", 16710 => "1110100100110010", 16711 => "0110111111001011", 16712 => "0110110101101011", 16713 => "0001101111001100", 16714 => "0001101100010110", 16715 => "0000000010110111", 16716 => "0101111001001000", 16717 => "1010010010100000", 16718 => "0111011011010110", 16719 => "1011001110001101", 16720 => "1110111010100100", 16721 => "0101001111111101", 16722 => "0100100010001000", 16723 => "1001011000010001", 16724 => "0011110100010100", 16725 => "1110000001100110", 16726 => "1101100010000000", 16727 => "0011010011011011", 16728 => "0001001001010101", 16729 => "0101110100111110", 16730 => "1000001010011000", 16731 => "1110110000100111", 16732 => "0011111101110010", 16733 => "0100001000111110", 16734 => "1100100011110011", 16735 => "1000011101010101", 16736 => "0011110011001010", 16737 => "1101110110010010", 16738 => "0111000101100100", 16739 => "0110110111000100", 16740 => "0111111000000100", 16741 => "0110001100101101", 16742 => "0110100111001101", 16743 => "1111010010110111", 16744 => "0001110001110110", 16745 => "1111110010100000", 16746 => "1011111101101011", 16747 => "0000011011010100", 16748 => "1100000011110011", 16749 => "0001110000010100", 16750 => "0100100001010111", 16751 => "1010001110010010", 16752 => "0101010000110001", 16753 => "1101100110011000", 16754 => "0110001111000110", 16755 => "0010100010011001", 16756 => "0100000001100001", 16757 => "0100101110110000", 16758 => "1001110101110100", 16759 => "0011011100011000", 16760 => "1101010101010101", 16761 => "1001011100100000", 16762 => "1010100001001101", 16763 => "0101100011110010", 16764 => "0111010110101010", 16765 => "1010101000001100", 16766 => "1010000001111100", 16767 => "1101100001111110", 16768 => "1111011000000011", 16769 => "0111111010011000", 16770 => "1111010100011011", 16771 => "0111001100101111", 16772 => "0101111001100100", 16773 => "1010001100111011", 16774 => "0100011110110111", 16775 => "0100011001011000", 16776 => "1111010000110001", 16777 => "1001110111101001", 16778 => "1100011100010111", 16779 => "0111101100000010", 16780 => "1000100110001100", 16781 => "0010001010111010", 16782 => "0111111001001100", 16783 => "0111110100110110", 16784 => "0101010010100011", 16785 => "0101110010100001", 16786 => "1000000111101011", 16787 => "0111101000110001", 16788 => "1001011111101110", 16789 => "0110000110010000", 16790 => "0101000000000010", 16791 => "1111010110000100", 16792 => "0101011110111111", 16793 => "0110000111011110", 16794 => "0000011101101010", 16795 => "0101011001001110", 16796 => "0000111101101010", 16797 => "0111111111010111", 16798 => "0100010101110001", 16799 => "1111001110011110", 16800 => "0001001110001101", 16801 => "1000111000111110", 16802 => "1110011001010111", 16803 => "0100111110101111", 16804 => "1100010010001001", 16805 => "1101000111010100", 16806 => "1001111111100110", 16807 => "0100000000001000", 16808 => "0000010100100110", 16809 => "0001001100010110", 16810 => "1000110101111010", 16811 => "1010001111101000", 16812 => "0110101000011110", 16813 => "0111110100001011", 16814 => "1110101001000001", 16815 => "0110011001110111", 16816 => "0001010111100011", 16817 => "1101111101100111", 16818 => "0100101100111111", 16819 => "1010111100000111", 16820 => "1111010010010011", 16821 => "0011010110100100", 16822 => "0110110011001010", 16823 => "1111100010001001", 16824 => "1011001011110101", 16825 => "1011110110110101", 16826 => "0101110101010010", 16827 => "1001111101100000", 16828 => "1111110001110001", 16829 => "1010101110110010", 16830 => "1010010011100011", 16831 => "1111001010100101", 16832 => "0101111001111000", 16833 => "0110100011100110", 16834 => "0100000011010010", 16835 => "0011100110011101", 16836 => "0000110010000011", 16837 => "0011100010011111", 16838 => "0100010011110001", 16839 => "0111100100011000", 16840 => "1010001111010001", 16841 => "1000010000010110", 16842 => "1101001001010000", 16843 => "1110110110011011", 16844 => "1001101011101010", 16845 => "0000000110100101", 16846 => "1110100000000010", 16847 => "0010110011110001", 16848 => "1111011000010010", 16849 => "1110100111001111", 16850 => "1011100010011010", 16851 => "1101011000011010", 16852 => "0100111000110111", 16853 => "1110110100010101", 16854 => "1001101110100101", 16855 => "0011111010101110", 16856 => "1010110011111110", 16857 => "1110101001101001", 16858 => "0010010100100110", 16859 => "1100100110011111", 16860 => "0010001100110011", 16861 => "1111000001000101", 16862 => "0000100111000111", 16863 => "0111000110000100", 16864 => "0111101110110011", 16865 => "0010111011011000", 16866 => "1010100111101101", 16867 => "0101101001001000", 16868 => "0101000101011011", 16869 => "0100111001110011", 16870 => "1001011000000011", 16871 => "0011010101100110", 16872 => "0110100110111110", 16873 => "0010111010001011", 16874 => "1010101000110000", 16875 => "0111000001111000", 16876 => "1101011110100010", 16877 => "0011000110001011", 16878 => "1000000001111000", 16879 => "0001110100011101", 16880 => "1001100010111001", 16881 => "1100100110101101", 16882 => "0011101111000111", 16883 => "0101001010110000", 16884 => "1010011011101101", 16885 => "0010011011110101", 16886 => "1011000101011111", 16887 => "1001010010001101", 16888 => "1000110111000001", 16889 => "1111001101100011", 16890 => "1000111101111001", 16891 => "0001010011110011", 16892 => "0011010101100101", 16893 => "0111010011110100", 16894 => "0011110111100000", 16895 => "0111101010011100", 16896 => "1011110101011110", 16897 => "0111001101010100", 16898 => "1100100100101010", 16899 => "1101010010111100", 16900 => "0100110001010111", 16901 => "1011000111111101", 16902 => "1100010010110111", 16903 => "1001001001100101", 16904 => "1111101001010011", 16905 => "1011111010100001", 16906 => "0010001111110001", 16907 => "0001010101110111", 16908 => "0101001010001010", 16909 => "1111000100111010", 16910 => "1010001111000001", 16911 => "1110000010111110", 16912 => "1101111001011001", 16913 => "0110011010011000", 16914 => "1001101000011110", 16915 => "1110100101101001", 16916 => "0110111101000001", 16917 => "0001000110111100", 16918 => "0101110111011101", 16919 => "0011010011001001", 16920 => "1101010110111111", 16921 => "0100100100101010", 16922 => "0100100110101111", 16923 => "0010100011111001", 16924 => "1100100010000101", 16925 => "1101000111101001", 16926 => "1100001100001011", 16927 => "1010111011011001", 16928 => "0111001101000101", 16929 => "1001111111000000", 16930 => "0010111100010011", 16931 => "1010000011101100", 16932 => "0001000110110100", 16933 => "1000100111001101", 16934 => "0100011101110101", 16935 => "0110111111111001", 16936 => "0100001101000111", 16937 => "1011111100111111", 16938 => "0111100011010000", 16939 => "0100101001001010", 16940 => "1101111100100001", 16941 => "1111011101110111", 16942 => "1100000101101111", 16943 => "0000111001011111", 16944 => "0000111000111000", 16945 => "0110001011000111", 16946 => "0001000111110000", 16947 => "1110100111001000", 16948 => "1110001010110000", 16949 => "1000000010100110", 16950 => "1000010011000101", 16951 => "0111011001110000", 16952 => "0001011101100011", 16953 => "0011100001110000", 16954 => "1011111110000111", 16955 => "0111010010000111", 16956 => "0011000101110000", 16957 => "1010110110001110", 16958 => "1000010010010000", 16959 => "1010101000011100", 16960 => "0000001100011110", 16961 => "1001010100011111", 16962 => "1100111000111110", 16963 => "0001100010101100", 16964 => "0001010011000110", 16965 => "0000000111001010", 16966 => "1000111100010001", 16967 => "1010111101011011", 16968 => "1001000011000100", 16969 => "0101000101111001", 16970 => "1001000001110010", 16971 => "1111001000110000", 16972 => "0011011001011010", 16973 => "0101100101011001", 16974 => "0110111010001001", 16975 => "1100001001110111", 16976 => "1011001010100011", 16977 => "1100110100001101", 16978 => "1111101110000010", 16979 => "1001011010110101", 16980 => "0101000110011101", 16981 => "1110001010011110", 16982 => "1111010111101100", 16983 => "1100000110100101", 16984 => "1001111011010110", 16985 => "1001010000111100", 16986 => "0000100110011000", 16987 => "0010001001010100", 16988 => "1011101111110001", 16989 => "1100011110111100", 16990 => "0111100011100010", 16991 => "1011111110111000", 16992 => "0110110100101000", 16993 => "0101100010111101", 16994 => "1011001011110110", 16995 => "0100101110100010", 16996 => "0000110111001100", 16997 => "1000101000000010", 16998 => "0000100110001010", 16999 => "0111000111001000", 17000 => "0111111001011001", 17001 => "0101001011111010", 17002 => "1110001110011111", 17003 => "1011000101100110", 17004 => "1010010110100101", 17005 => "0111110101010111", 17006 => "1111101111001101", 17007 => "0110011000010101", 17008 => "1011010100100001", 17009 => "1111100101000100", 17010 => "1001110001100111", 17011 => "0110010101110010", 17012 => "0111010100110111", 17013 => "1110001010101011", 17014 => "1011011010110100", 17015 => "0011110011101100", 17016 => "0001011001100010", 17017 => "0101110000010111", 17018 => "1111101101111010", 17019 => "0000111100101111", 17020 => "0111011010001011", 17021 => "1110110011000001", 17022 => "0100101111101010", 17023 => "1010000001111100", 17024 => "1100010001110001", 17025 => "0011001111110101", 17026 => "0111111000100001", 17027 => "0101011100011101", 17028 => "1110111000001001", 17029 => "0110000010011110", 17030 => "1111110000010010", 17031 => "0101000101111000", 17032 => "0000011011011111", 17033 => "1000100100001000", 17034 => "1011110101011100", 17035 => "0010110111101011", 17036 => "1000001011100111", 17037 => "1111000000010100", 17038 => "0011010010100010", 17039 => "1100100111011001", 17040 => "0110101110111000", 17041 => "0100100111001001", 17042 => "1000110010011010", 17043 => "0000100110111100", 17044 => "1101110110101101", 17045 => "0110010001001010", 17046 => "0010111111100001", 17047 => "0011011100111010", 17048 => "0111001010110111", 17049 => "1110111011111111", 17050 => "0101000011000001", 17051 => "1000011111101011", 17052 => "1011000100111111", 17053 => "1111111001011011", 17054 => "0111111111011111", 17055 => "0001011100010011", 17056 => "1111110111000010", 17057 => "0110111110011100", 17058 => "1101000010011111", 17059 => "0011111011101010", 17060 => "1111111010001110", 17061 => "0101101101011110", 17062 => "0000101001011010", 17063 => "1010100000000101", 17064 => "0110101011000010", 17065 => "0000111100110111", 17066 => "1000000100101000", 17067 => "1011110101000000", 17068 => "0111100111011011", 17069 => "1110111000000000", 17070 => "1110011000111000", 17071 => "0010101010111001", 17072 => "1000001001001001", 17073 => "0011001001111011", 17074 => "1011101001111111", 17075 => "0011111000110000", 17076 => "1001000000010111", 17077 => "0001101000100000", 17078 => "0101010010100001", 17079 => "1111111101000000", 17080 => "0110011010101110", 17081 => "0101110111110010", 17082 => "0110000011010111", 17083 => "1101011000111010", 17084 => "1111001100111010", 17085 => "1011011001011110", 17086 => "0101011101100000", 17087 => "1101111110011011", 17088 => "0100110000101101", 17089 => "0001100100011001", 17090 => "1100100000000000", 17091 => "1010100001000000", 17092 => "0000010111001101", 17093 => "0011101010110010", 17094 => "1000110011101001", 17095 => "0000110110000110", 17096 => "0110010111111101", 17097 => "1110000100111110", 17098 => "1010010010010110", 17099 => "0011111000110001", 17100 => "1000101010001011", 17101 => "1010100011010001", 17102 => "0101111111001011", 17103 => "1000110001100010", 17104 => "0100111000101101", 17105 => "0011101110110100", 17106 => "1101110010011000", 17107 => "0000001010100001", 17108 => "0011011001011000", 17109 => "1110000100010001", 17110 => "1101010000010111", 17111 => "0010111100110001", 17112 => "0100011100100101", 17113 => "0111000001010010", 17114 => "1000001101010100", 17115 => "1111010001110011", 17116 => "0000100010000110", 17117 => "1110110000001000", 17118 => "1110110000001010", 17119 => "0101011111010001", 17120 => "1100110001000110", 17121 => "0111000111001000", 17122 => "1010101110101111", 17123 => "0010101101110111", 17124 => "1101001010010110", 17125 => "0000011100111101", 17126 => "1100111010010101", 17127 => "1011000100010100", 17128 => "1110001000110111", 17129 => "1010000011010010", 17130 => "0101110110001101", 17131 => "1111110011011111", 17132 => "1011110001100110", 17133 => "1101000011110100", 17134 => "1101000000100010", 17135 => "0101111000101001", 17136 => "1000110101001001", 17137 => "1001101101111011", 17138 => "0110111000001000", 17139 => "1000000101101010", 17140 => "1100000100111011", 17141 => "1110001001000011", 17142 => "1101110111100101", 17143 => "0001010100110101", 17144 => "1110010010100100", 17145 => "1101101100101010", 17146 => "0010010010010100", 17147 => "1011111010110101", 17148 => "1010100101011000", 17149 => "1111000011111110", 17150 => "1001001000110100", 17151 => "1010010101110000", 17152 => "1011010100000000", 17153 => "0101101010001010", 17154 => "0111011001111000", 17155 => "0010001101111111", 17156 => "0001111111001011", 17157 => "1111100111010011", 17158 => "1111010100001000", 17159 => "0110010110110111", 17160 => "0001110100010100", 17161 => "0010010010010010", 17162 => "1011010110100010", 17163 => "1001010001111110", 17164 => "1001000011000101", 17165 => "0000010101010000", 17166 => "0000000110011100", 17167 => "1110000000001110", 17168 => "0111010000101010", 17169 => "0110001111011111", 17170 => "1110010101110010", 17171 => "1110110011100100", 17172 => "0111011111111000", 17173 => "1101000010111000", 17174 => "0111000010000000", 17175 => "0101101110000101", 17176 => "1001111111111101", 17177 => "1011111011000110", 17178 => "0011101010110110", 17179 => "1110000000101011", 17180 => "0100000101010010", 17181 => "1111010000111011", 17182 => "0001101011010100", 17183 => "0110010011010100", 17184 => "0100101101101101", 17185 => "0011000001101010", 17186 => "0010111000010110", 17187 => "0100010011011000", 17188 => "1000000100110001", 17189 => "0111011110111001", 17190 => "0011001010111100", 17191 => "0010011000000110", 17192 => "1110100000111110", 17193 => "0100111010010101", 17194 => "0111011100011110", 17195 => "1100101000010011", 17196 => "1001110111111011", 17197 => "1111001010000110", 17198 => "0111001010101010", 17199 => "0111111111001110", 17200 => "1000000000011010", 17201 => "0001100101000010", 17202 => "1111101111111101", 17203 => "0000110111110010", 17204 => "1011010111010110", 17205 => "0010001101011001", 17206 => "1001001111001101", 17207 => "1111111000010011", 17208 => "0101111010101100", 17209 => "0001110001001010", 17210 => "0111010101011101", 17211 => "1001100001101011", 17212 => "1010111100000110", 17213 => "0111000111010011", 17214 => "1000100110100011", 17215 => "0010111110011000", 17216 => "0000111110111000", 17217 => "1000010000110000", 17218 => "1001110111111110", 17219 => "0111011101111010", 17220 => "0111100011101100", 17221 => "0001101100011100", 17222 => "1010011101011000", 17223 => "0000111100011001", 17224 => "1011010000101101", 17225 => "0101000100100110", 17226 => "0111111000100101", 17227 => "1001101100101001", 17228 => "0111111001000011", 17229 => "1001011000100010", 17230 => "0100100010011100", 17231 => "0011010011110111", 17232 => "1010110100100101", 17233 => "1011001110000100", 17234 => "0110010011101000", 17235 => "0100001011001000", 17236 => "1110010101110111", 17237 => "1111100101000101", 17238 => "0101100101110100", 17239 => "0000011110010011", 17240 => "0001110100111011", 17241 => "1111111100011000", 17242 => "1000000110110000", 17243 => "1111001000000001", 17244 => "0111000111011000", 17245 => "0001111011111101", 17246 => "0000010000111100", 17247 => "0000011000100010", 17248 => "1010000001000001", 17249 => "0110001010101000", 17250 => "0101111101100110", 17251 => "1011111101110110", 17252 => "1011010111100100", 17253 => "1010101011001111", 17254 => "0111110100110111", 17255 => "1111001100101001", 17256 => "1000011011100001", 17257 => "0100101111100101", 17258 => "1001001110000110", 17259 => "0101001111000111", 17260 => "1011110100101110", 17261 => "0000001111000000", 17262 => "0101110100101111", 17263 => "1000001101001110", 17264 => "0111110001011100", 17265 => "1100101011010110", 17266 => "0000111011111101", 17267 => "0000111110100101", 17268 => "0100101100101010", 17269 => "0111100001100110", 17270 => "1000010000100000", 17271 => "1000110000010001", 17272 => "1110111011000001", 17273 => "0000000001000010", 17274 => "1001100000011011", 17275 => "1100000110000111", 17276 => "1100101001000000", 17277 => "1001101101100000", 17278 => "0111110101100000", 17279 => "1110111101110110", 17280 => "1010011100111011", 17281 => "0010011011110010", 17282 => "1011100000000110", 17283 => "1101111011000001", 17284 => "1010001100001101", 17285 => "1011001111010111", 17286 => "1111101001110010", 17287 => "0100111000110010", 17288 => "1010100011111111", 17289 => "1110111011000001", 17290 => "0011001101011110", 17291 => "0111000010000110", 17292 => "1111001000100101", 17293 => "1101110100100010", 17294 => "1111001100100110", 17295 => "0011110100100010", 17296 => "1111011111011100", 17297 => "0001010111100011", 17298 => "0111001011101111", 17299 => "1000011111101111", 17300 => "0101000101000001", 17301 => "0010111001101110", 17302 => "0001110110111111", 17303 => "1100100011011110", 17304 => "0100100000100001", 17305 => "0000110111010100", 17306 => "1101001110111111", 17307 => "1001111101110110", 17308 => "1111111111001010", 17309 => "0010111111001111", 17310 => "1100101010000100", 17311 => "1100001000011010", 17312 => "0111001110100111", 17313 => "0101110111101111", 17314 => "1100011101100011", 17315 => "0101100000000011", 17316 => "1110101101100000", 17317 => "0111001110010100", 17318 => "1100110100101000", 17319 => "1100001000110011", 17320 => "1110101111000110", 17321 => "0000101000001001", 17322 => "0001001010001001", 17323 => "0001110100110011", 17324 => "0011001001011000", 17325 => "1110101111011011", 17326 => "1011110110001100", 17327 => "1001110011011000", 17328 => "1111011110100111", 17329 => "0000100111011010", 17330 => "1001010010101011", 17331 => "0100100011000100", 17332 => "0111101100000000", 17333 => "0101001000110110", 17334 => "0101001000010001", 17335 => "1000100010100011", 17336 => "1000000110110101", 17337 => "0011101001110111", 17338 => "1111000100100001", 17339 => "0001100111101110", 17340 => "1110100001001101", 17341 => "0010000111000000", 17342 => "1101100000100110", 17343 => "0010101001100011", 17344 => "0001011010110001", 17345 => "1101001110000001", 17346 => "0000111000001001", 17347 => "1100110101000001", 17348 => "1000001100000101", 17349 => "1101110111111000", 17350 => "0101010000011001", 17351 => "1000010001001100", 17352 => "1010100010001111", 17353 => "1001011000011001", 17354 => "0110010101000111", 17355 => "1000100110110011", 17356 => "1010101011101000", 17357 => "0111011100100001", 17358 => "1100001000110010", 17359 => "1101010010110100", 17360 => "1101110011101100", 17361 => "0110111111000100", 17362 => "0101000101101001", 17363 => "1111100101010010", 17364 => "1011010111001011", 17365 => "1101000101001001", 17366 => "1100111000000101", 17367 => "0110011010000001", 17368 => "1011001000111010", 17369 => "1011110101101011", 17370 => "1000100100011010", 17371 => "0111111000011001", 17372 => "1011001011100110", 17373 => "0001110011100101", 17374 => "0110001100010110", 17375 => "0110001100000110", 17376 => "0100011010101101", 17377 => "1101100010110111", 17378 => "1110101011001010", 17379 => "1000011111011110", 17380 => "1011111010000000", 17381 => "0010110111010001", 17382 => "0010001000101001", 17383 => "1110111101101000", 17384 => "0111101011001001", 17385 => "1110110110001111", 17386 => "1001110101100000", 17387 => "1011111001010100", 17388 => "1011011101100111", 17389 => "0000010010000100", 17390 => "0000000000000000", 17391 => "1011100111001010", 17392 => "1011111100001101", 17393 => "1111110110101110", 17394 => "1110001101000111", 17395 => "1001100110110001", 17396 => "1110010000101111", 17397 => "1001111111001000", 17398 => "0011010111001101", 17399 => "0010100100001101", 17400 => "0000010000100011", 17401 => "1101010101111111", 17402 => "1111100010101001", 17403 => "1010111111010001", 17404 => "0100101100110101", 17405 => "0110101001100010", 17406 => "0010110010101010", 17407 => "0101100000110110", 17408 => "0110100111010100", 17409 => "0111010001111111", 17410 => "0001001010000011", 17411 => "0001010101111010", 17412 => "0111110100100001", 17413 => "0110001010101011", 17414 => "1111001110010011", 17415 => "1011111110000111", 17416 => "0101101010010000", 17417 => "1100010111011101", 17418 => "1111110011000110", 17419 => "0011111010110011", 17420 => "1011111010010010", 17421 => "0010011001111110", 17422 => "1010111000100111", 17423 => "1101010000111010", 17424 => "1100000111000111", 17425 => "0110111100000000", 17426 => "1110001011111110", 17427 => "0001000010101011", 17428 => "0111100111101100", 17429 => "1000010010101011", 17430 => "1111010000101100", 17431 => "1110010011001000", 17432 => "0010000010010011", 17433 => "1001110111000110", 17434 => "1010100000111100", 17435 => "1110011111010101", 17436 => "1000011100011100", 17437 => "0010001101101010", 17438 => "0010110111111111", 17439 => "0000111001001001", 17440 => "1101111101000000", 17441 => "0010000000001010", 17442 => "0110010011111010", 17443 => "1111001001000000", 17444 => "0011000101110010", 17445 => "0010010110101010", 17446 => "0000011100100100", 17447 => "1001000111110001", 17448 => "1000110011111110", 17449 => "1110000011101001", 17450 => "1010011011100101", 17451 => "0100110001011010", 17452 => "0111101111111100", 17453 => "0110010100011001", 17454 => "1011010001001010", 17455 => "1010010001110100", 17456 => "1010110001101001", 17457 => "0000100000001001", 17458 => "1011100101111111", 17459 => "1110111000011110", 17460 => "0101100001100010", 17461 => "1010101111110110", 17462 => "0001101100000100", 17463 => "1111111110110011", 17464 => "0101000010000001", 17465 => "1101011101111001", 17466 => "0001101111111110", 17467 => "1000101101011000", 17468 => "0110110011000110", 17469 => "1011010011111110", 17470 => "0010000001000110", 17471 => "0101011100010001", 17472 => "0101011000000000", 17473 => "0000001111111101", 17474 => "1111000111101001", 17475 => "1000001111111101", 17476 => "0011101001111011", 17477 => "0010101101100011", 17478 => "0011011111001101", 17479 => "1001110010000011", 17480 => "1010011111000011", 17481 => "1010000101100110", 17482 => "1100001110100101", 17483 => "1100001111110110", 17484 => "1100001011101111", 17485 => "1101011110100000", 17486 => "1101110001111111", 17487 => "0011010001010101", 17488 => "0100100011000110", 17489 => "1000001001011110", 17490 => "0110110000010011", 17491 => "1001100001000011", 17492 => "0100111100001010", 17493 => "1001100011010010", 17494 => "1110100101010110", 17495 => "0110011010011001", 17496 => "1010110011101001", 17497 => "0111100100001000", 17498 => "1101110111101011", 17499 => "0111010100101111", 17500 => "1111001010110100", 17501 => "1001001100100010", 17502 => "1010100001110100", 17503 => "0001110111011000", 17504 => "0100010001110110", 17505 => "0100100010100101", 17506 => "1101001001010011", 17507 => "1010010000001101", 17508 => "0011110000011101", 17509 => "1100001111001000", 17510 => "0011001111100110", 17511 => "0010111001001010", 17512 => "0110011001000000", 17513 => "1001111010010000", 17514 => "1000010001011110", 17515 => "1101011001001101", 17516 => "1101010000111101", 17517 => "0101001011010011", 17518 => "0011111000111000", 17519 => "1010101010101001", 17520 => "0111010011010011", 17521 => "0001100111100000", 17522 => "1101100001011001", 17523 => "0100010010110110", 17524 => "0000011011101111", 17525 => "0010010010010000", 17526 => "1101011011101011", 17527 => "0100010111011100", 17528 => "0001001100011001", 17529 => "1100100001110000", 17530 => "0100010011010101", 17531 => "0011111111010101", 17532 => "0111101110010011", 17533 => "0101111010011111", 17534 => "0100101100010100", 17535 => "1000111011110111", 17536 => "1100000100010010", 17537 => "1110111101111011", 17538 => "0010010111010010", 17539 => "1011110000001110", 17540 => "0110010010110010", 17541 => "0111110111111010", 17542 => "0111110100001000", 17543 => "0111100111010111", 17544 => "1110010010110011", 17545 => "1011011111011010", 17546 => "0000110011111100", 17547 => "0110111100011100", 17548 => "0011011110010110", 17549 => "1110001000100011", 17550 => "0100010010011000", 17551 => "0111011111101101", 17552 => "1101011110000001", 17553 => "1111110111111010", 17554 => "0011010100000101", 17555 => "0010010100111110", 17556 => "0110101101010111", 17557 => "0111001110110110", 17558 => "1011111000010001", 17559 => "1100101001111111", 17560 => "1000001011011100", 17561 => "1001000001110111", 17562 => "1111101101010110", 17563 => "0111111110001010", 17564 => "1111110011101001", 17565 => "1101010001011000", 17566 => "1101000101001100", 17567 => "0101001110101110", 17568 => "0100001011000111", 17569 => "0000111110011000", 17570 => "1100001000011000", 17571 => "1100110101101101", 17572 => "1111100000110100", 17573 => "0011010011100100", 17574 => "1111011000010100", 17575 => "0101110100111110", 17576 => "1000101001011111", 17577 => "0011000101110111", 17578 => "1010111111000001", 17579 => "1110001001001100", 17580 => "0000010010000001", 17581 => "0111000011000011", 17582 => "1011101000101101", 17583 => "1000110001111100", 17584 => "0000011000001001", 17585 => "0111010111011110", 17586 => "0111100011010011", 17587 => "1000100001011011", 17588 => "1001010111001011", 17589 => "1111101110001111", 17590 => "0011110100001111", 17591 => "1000010001111100", 17592 => "0001100000100111", 17593 => "0010110111111000", 17594 => "1111110011010110", 17595 => "0010000111111001", 17596 => "0110001101110110", 17597 => "1110010100011110", 17598 => "1100111110000010", 17599 => "1101001010100000", 17600 => "1111000010100110", 17601 => "0111001100100111", 17602 => "0001000101110011", 17603 => "0010011011010110", 17604 => "0000000010101000", 17605 => "0000111011111001", 17606 => "0100000010111010", 17607 => "1000000011101101", 17608 => "0110110001100011", 17609 => "1000011011000110", 17610 => "1011101001010010", 17611 => "0110111100011010", 17612 => "1100000000100010", 17613 => "1001111001000001", 17614 => "1111100101010101", 17615 => "1001000101001010", 17616 => "1110101010010111", 17617 => "0000111101000010", 17618 => "1111100000100010", 17619 => "1111110111110010", 17620 => "1110101111100011", 17621 => "0101010101101000", 17622 => "1000011010111011", 17623 => "0111001011111011", 17624 => "0110000110110100", 17625 => "0011101001110100", 17626 => "1001001000001100", 17627 => "0100001111101111", 17628 => "1001011001111101", 17629 => "0000110110011011", 17630 => "1110010010100011", 17631 => "0010101001110001", 17632 => "0001111111110100", 17633 => "0010000000010100", 17634 => "0111110101000111", 17635 => "0011000111110101", 17636 => "0011100110100111", 17637 => "1100001101111101", 17638 => "1111010100111010", 17639 => "0001011111000111", 17640 => "1011010111000100", 17641 => "1111110110001111", 17642 => "1001100110101011", 17643 => "1001010110111000", 17644 => "1111001110110000", 17645 => "0110101000010001", 17646 => "1101011000100011", 17647 => "1100001110001001", 17648 => "1000101111101000", 17649 => "0000010010000011", 17650 => "0010101110100101", 17651 => "0010001100100100", 17652 => "1111010100011000", 17653 => "0010001101001101", 17654 => "1001101110100100", 17655 => "0000110001000111", 17656 => "1101100000100110", 17657 => "1011010111101000", 17658 => "1000001100100000", 17659 => "1110111011001001", 17660 => "0100001110011111", 17661 => "0110010111010100", 17662 => "0111011111100000", 17663 => "1110100010100011", 17664 => "0100011111100001", 17665 => "0110101101110000", 17666 => "1011100010110001", 17667 => "1111010110001110", 17668 => "1000000100110001", 17669 => "1100000101100011", 17670 => "1111000011101001", 17671 => "1001101110011001", 17672 => "0100111010000100", 17673 => "1010101011010110", 17674 => "0011010110111101", 17675 => "1101001001011011", 17676 => "0111000101001010", 17677 => "1111000000110100", 17678 => "0110101011000101", 17679 => "0000111001011100", 17680 => "1010100000010011", 17681 => "1001100100010111", 17682 => "1100010001100000", 17683 => "0100001101011010", 17684 => "1011001101101110", 17685 => "1111100111011100", 17686 => "1111110111110000", 17687 => "1110110100011100", 17688 => "0110101011101000", 17689 => "1100010010111011", 17690 => "0110101000010101", 17691 => "1111011011100001", 17692 => "0001000011100110", 17693 => "0110010010100111", 17694 => "1100110001110110", 17695 => "1001100111010001", 17696 => "1100011101100100", 17697 => "0100100110100010", 17698 => "1110011000010001", 17699 => "0011001000001100", 17700 => "1101010000000010", 17701 => "0111111101101101", 17702 => "1100110100010110", 17703 => "1110011101111001", 17704 => "1100010001001010", 17705 => "1010111101110001", 17706 => "1010101111100011", 17707 => "0000101010011000", 17708 => "0110010011110000", 17709 => "0100000100100011", 17710 => "1010010000000001", 17711 => "1100001100011000", 17712 => "0000010110001100", 17713 => "0000011111011011", 17714 => "0100111011001110", 17715 => "1100110011000110", 17716 => "0011100111000101", 17717 => "1010110010010100", 17718 => "0001010000100000", 17719 => "1011100111101010", 17720 => "1111111111100100", 17721 => "1000011011100111", 17722 => "0100101101011101", 17723 => "0111000010110111", 17724 => "1000111101011001", 17725 => "1110001101001010", 17726 => "0100100000011110", 17727 => "0100111000110100", 17728 => "0000100000111100", 17729 => "1000011101111010", 17730 => "1001101010111011", 17731 => "1010101101001101", 17732 => "0010010001100001", 17733 => "0010111010000010", 17734 => "1001000100100110", 17735 => "0100100000101000", 17736 => "0000011110011111", 17737 => "1000100111100001", 17738 => "1111111001010000", 17739 => "0110010010010111", 17740 => "0001100010000101", 17741 => "1011111100010101", 17742 => "1010111111111101", 17743 => "0000010101111110", 17744 => "1101110000100001", 17745 => "1000000111010111", 17746 => "1101010010111111", 17747 => "0110010001100100", 17748 => "0110111110000111", 17749 => "1010100011001101", 17750 => "0101011101011111", 17751 => "0111001001110110", 17752 => "0111011000000110", 17753 => "1111111100110010", 17754 => "1110101001101101", 17755 => "1111100010010101", 17756 => "0011101000001111", 17757 => "0001000010011110", 17758 => "1011000110011010", 17759 => "1101010001011100", 17760 => "0001100100010101", 17761 => "1111110101011110", 17762 => "1001001011000101", 17763 => "1010110011110110", 17764 => "0100000110110110", 17765 => "1111101111000111", 17766 => "0011100111010011", 17767 => "1101100001000010", 17768 => "0010111101010001", 17769 => "0001001101000100", 17770 => "0110110100011101", 17771 => "1010001000001001", 17772 => "0110111100101100", 17773 => "0110000101000000", 17774 => "0110110111100001", 17775 => "1010110110001011", 17776 => "0001011000000011", 17777 => "0010010011001000", 17778 => "0111110111001101", 17779 => "1110100101011101", 17780 => "1111000000000010", 17781 => "1111001111011001", 17782 => "0110000010110100", 17783 => "0110101011010110", 17784 => "1001001010001010", 17785 => "0111010011110100", 17786 => "0011011011100100", 17787 => "1010001001000010", 17788 => "1000110011000011", 17789 => "0010111101000011", 17790 => "1111010010100010", 17791 => "1101011101111101", 17792 => "0011001110111111", 17793 => "0010101000000101", 17794 => "0110100111001011", 17795 => "1110000110010010", 17796 => "0010111100001100", 17797 => "0100111010001111", 17798 => "0101101010010010", 17799 => "1110110001001101", 17800 => "0110110101100101", 17801 => "0011011001111001", 17802 => "1111100110001010", 17803 => "1001100000100101", 17804 => "1100101110111010", 17805 => "1100111010110000", 17806 => "0101001110101111", 17807 => "1101110000010001", 17808 => "0011011110111111", 17809 => "1110010001110110", 17810 => "0111000101111010", 17811 => "0011001010000110", 17812 => "1011010111010100", 17813 => "0100111011010001", 17814 => "1010011110100101", 17815 => "0110000111011111", 17816 => "1001111110000000", 17817 => "1010111110010010", 17818 => "0110011011101011", 17819 => "1100100110000110", 17820 => "0110000101011110", 17821 => "1010010111100110", 17822 => "1101011000010001", 17823 => "1001011001000101", 17824 => "1110111111000110", 17825 => "1011100100100010", 17826 => "0111111011100000", 17827 => "0011000001101111", 17828 => "0101110001011011", 17829 => "1001001100000001", 17830 => "1111100001001000", 17831 => "1101011001111101", 17832 => "0110100110101001", 17833 => "0011010000001011", 17834 => "0001010000101000", 17835 => "1101100001010101", 17836 => "1001000001001010", 17837 => "1100110010001111", 17838 => "0101000111100100", 17839 => "0011001111110101", 17840 => "0011110111101001", 17841 => "0011001001001110", 17842 => "1011101110100001", 17843 => "0101110010111101", 17844 => "1101010000100110", 17845 => "1110000010100010", 17846 => "0100101000111011", 17847 => "0100111101101000", 17848 => "1101000010000000", 17849 => "1010101101010110", 17850 => "0110110111010111", 17851 => "1010011001011101", 17852 => "1110000110100000", 17853 => "0000010001000011", 17854 => "0010010100011101", 17855 => "1011000101111000", 17856 => "1000110010100011", 17857 => "1001001111110110", 17858 => "0101110101110100", 17859 => "0011111111001011", 17860 => "1000000011000101", 17861 => "0111000101000111", 17862 => "1100110110010000", 17863 => "0110000010011010", 17864 => "0010010001101111", 17865 => "0011001010000110", 17866 => "0001011001001111", 17867 => "0101010001010101", 17868 => "0001000110100011", 17869 => "1111100111100001", 17870 => "1110100010001100", 17871 => "0111011100101000", 17872 => "0101110010001011", 17873 => "0111100110110110", 17874 => "1011101000010011", 17875 => "1000110110101011", 17876 => "0000110101101101", 17877 => "1010011001001100", 17878 => "0101001101011011", 17879 => "0100101001001110", 17880 => "1110110100000000", 17881 => "0110111011011011", 17882 => "0100011111111100", 17883 => "0000010110000110", 17884 => "0000010111100110", 17885 => "0111010010100101", 17886 => "1110000100110101", 17887 => "0100100000111010", 17888 => "0101100000100000", 17889 => "0010101100111111", 17890 => "1000011010011111", 17891 => "0000001000001101", 17892 => "1100000101001111", 17893 => "1111101101011000", 17894 => "1101110111110110", 17895 => "1011011010001100", 17896 => "1011001011011100", 17897 => "0100011000000100", 17898 => "0001011011110010", 17899 => "0011100011101110", 17900 => "1000011111000000", 17901 => "1011110111111011", 17902 => "1000000100000111", 17903 => "0101110001000111", 17904 => "1100010000111111", 17905 => "1010101001011011", 17906 => "0111111001100101", 17907 => "1010100111100101", 17908 => "1010001000111001", 17909 => "1111100110100010", 17910 => "0000101010011101", 17911 => "0100111000101110", 17912 => "1011011000101010", 17913 => "0101011110111000", 17914 => "0101011111101010", 17915 => "1111100111010100", 17916 => "0100010000001101", 17917 => "0010111110000111", 17918 => "0111110111001101", 17919 => "0010011111011111", 17920 => "0011010100111101", 17921 => "0111001001111000", 17922 => "0011000111010001", 17923 => "1110101001100001", 17924 => "0000110000011001", 17925 => "0011001110010000", 17926 => "0111110101000001", 17927 => "1111111001111011", 17928 => "0100100100011010", 17929 => "1011100100001110", 17930 => "1111000010011111", 17931 => "1010000010000100", 17932 => "0001110011111010", 17933 => "1010011001100000", 17934 => "0011001011100010", 17935 => "0101000100011010", 17936 => "0100001001110000", 17937 => "1001011111101100", 17938 => "0010101001011010", 17939 => "0110100000100000", 17940 => "1011101011101100", 17941 => "0110101000111000", 17942 => "1101101000101110", 17943 => "1110100000010000", 17944 => "1011101001000101", 17945 => "1001101011111000", 17946 => "0100111100001000", 17947 => "1110001010110101", 17948 => "0110101011010100", 17949 => "0000101111001111", 17950 => "0011110111101000", 17951 => "1110111000111111", 17952 => "1110011100010111", 17953 => "0010100011111111", 17954 => "0100100001111111", 17955 => "0100100101010010", 17956 => "0000010010000000", 17957 => "1110110011000111", 17958 => "1111111010000010", 17959 => "1000001011101110", 17960 => "1001001100010010", 17961 => "0100111110100001", 17962 => "1111011110000011", 17963 => "0000000101011100", 17964 => "0001001000001110", 17965 => "1101111101010101", 17966 => "1101111101110000", 17967 => "1010010110100001", 17968 => "0010000010011011", 17969 => "0111101111010011", 17970 => "1010101011100011", 17971 => "1000111000010111", 17972 => "0111101100101010", 17973 => "1010110011001110", 17974 => "1000011010010110", 17975 => "0010111010100001", 17976 => "0111001001100100", 17977 => "1011100100001010", 17978 => "0100000110000001", 17979 => "1000100001110000", 17980 => "0010000111001010", 17981 => "0100111101010101", 17982 => "1011010100001111", 17983 => "1000100101011000", 17984 => "1101110011010010", 17985 => "1101000100000001", 17986 => "1110111001001111", 17987 => "0010010110110010", 17988 => "1100001001110110", 17989 => "0000101010010100", 17990 => "1101010101111011", 17991 => "1101001000001001", 17992 => "0100011101100011", 17993 => "1011011000100101", 17994 => "0100100101101101", 17995 => "1001101011101110", 17996 => "1001010110101100", 17997 => "0100010001101101", 17998 => "1100110000011010", 17999 => "0100010001111011", 18000 => "0010001111001111", 18001 => "1011111100100111", 18002 => "1111100010000110", 18003 => "1010010100110000", 18004 => "0111010101111111", 18005 => "1011001101011001", 18006 => "1111001100111011", 18007 => "1000000011010000", 18008 => "0011111001010101", 18009 => "1111100001100011", 18010 => "0011100101010111", 18011 => "1001100111110101", 18012 => "1100001110111101", 18013 => "1101010000110011", 18014 => "1101011110000011", 18015 => "1010010111100010", 18016 => "0111001110000101", 18017 => "0100010011110011", 18018 => "1001011110000110", 18019 => "0101001001101101", 18020 => "1110010100010000", 18021 => "0000101101111110", 18022 => "0101100101011110", 18023 => "0110010110001001", 18024 => "0110010001101011", 18025 => "1100100010110010", 18026 => "1010000010101010", 18027 => "1100111010101100", 18028 => "0011111010000110", 18029 => "1111001011001111", 18030 => "0111011011010110", 18031 => "0110001000001011", 18032 => "0100000100101010", 18033 => "1010010100100101", 18034 => "0010101100010110", 18035 => "1110001101100110", 18036 => "0010011111111001", 18037 => "0101001001011100", 18038 => "0001010101000110", 18039 => "0010110001111011", 18040 => "1110110010101010", 18041 => "1001011101000000", 18042 => "0001101100110001", 18043 => "0000011001010110", 18044 => "0001111101011000", 18045 => "0110100110110001", 18046 => "1101010011101011", 18047 => "1100110000101100", 18048 => "0001011111110001", 18049 => "0101001110001101", 18050 => "1001001110011001", 18051 => "1000101011111001", 18052 => "0000101101101011", 18053 => "0011100111100011", 18054 => "0111110110101010", 18055 => "0110100100101001", 18056 => "1110100000111100", 18057 => "0110100010010000", 18058 => "1100100101010101", 18059 => "0101010111101011", 18060 => "0110001101010011", 18061 => "0010101010110001", 18062 => "1001011101001111", 18063 => "1010110101111101", 18064 => "1100111110111110", 18065 => "1001100110011110", 18066 => "0011010011010110", 18067 => "0001101101111010", 18068 => "0110110111001110", 18069 => "0111001000101011", 18070 => "1000011010101000", 18071 => "1101000100100110", 18072 => "0011110010111101", 18073 => "0101001000100101", 18074 => "0111101001001000", 18075 => "0101001001000101", 18076 => "0011110011101001", 18077 => "0001010001110111", 18078 => "1100110000001001", 18079 => "0011111101011000", 18080 => "0001110011010011", 18081 => "1001111111001001", 18082 => "0010101000100001", 18083 => "0011010010011110", 18084 => "1110100000000110", 18085 => "1100111000111111", 18086 => "0110110001000011", 18087 => "1110101001011111", 18088 => "1110111111011100", 18089 => "0101001110111100", 18090 => "1000101001111110", 18091 => "0111100101111011", 18092 => "0111000100011101", 18093 => "0111110101111011", 18094 => "1010110100000001", 18095 => "1000010010010101", 18096 => "1011100110110010", 18097 => "0011100110110110", 18098 => "1100010000000111", 18099 => "1111011011000011", 18100 => "0011100110011011", 18101 => "1000101100011111", 18102 => "1011000010010000", 18103 => "0011101000110111", 18104 => "1101000001101110", 18105 => "0111001101110100", 18106 => "1010110100001001", 18107 => "1000100000110001", 18108 => "1101110110011111", 18109 => "1000011001100010", 18110 => "1001011111111011", 18111 => "1111000101010111", 18112 => "0111010001111011", 18113 => "0110000101011111", 18114 => "0110101000000111", 18115 => "0101100101111101", 18116 => "0010101110111010", 18117 => "1110100000001010", 18118 => "1000110011010001", 18119 => "1011011111100110", 18120 => "0010101000101111", 18121 => "0111110011001001", 18122 => "1010001100101000", 18123 => "1100000110111011", 18124 => "0010011111101111", 18125 => "0010101101000110", 18126 => "1001111000000011", 18127 => "0110100010011001", 18128 => "1001101010101000", 18129 => "0110010001101100", 18130 => "0100100001010111", 18131 => "1101110101000110", 18132 => "0110100111110100", 18133 => "1111001000111111", 18134 => "0110110111001000", 18135 => "0110001010000111", 18136 => "0100110101000101", 18137 => "1110001010001010", 18138 => "0110000101010011", 18139 => "1101010010111100", 18140 => "0110000001100010", 18141 => "1111110000110100", 18142 => "0101011101011011", 18143 => "0011001001010001", 18144 => "1010100110100001", 18145 => "0101110001011001", 18146 => "0001010100010100", 18147 => "0000110001011100", 18148 => "1110100000011001", 18149 => "1011110001101110", 18150 => "1100111010111001", 18151 => "1111010111110001", 18152 => "1001000101011001", 18153 => "1001111111111001", 18154 => "1101001110100000", 18155 => "1010111001100111", 18156 => "0101000110100010", 18157 => "1110111111010011", 18158 => "0101111010100100", 18159 => "0111110001000111", 18160 => "1000011111111101", 18161 => "0011001110110110", 18162 => "0100011101100100", 18163 => "1110011100011110", 18164 => "0010110100100111", 18165 => "0001111011000001", 18166 => "0111111000110111", 18167 => "0011010110100100", 18168 => "1110011000111011", 18169 => "0111010000100100", 18170 => "1010100000100100", 18171 => "0001001011100110", 18172 => "0100001001101111", 18173 => "1100001011101010", 18174 => "1100101011000011", 18175 => "1010011110010111", 18176 => "1010001101011100", 18177 => "1100011101101001", 18178 => "0110010110000001", 18179 => "0110111110100011", 18180 => "1111000111110101", 18181 => "0011101110101001", 18182 => "1111111010001011", 18183 => "0010100011001011", 18184 => "1011101001010101", 18185 => "1001101110011000", 18186 => "1000110111010001", 18187 => "0110111100011010", 18188 => "0100111011101011", 18189 => "1110000001001101", 18190 => "1100100110001111", 18191 => "0110101111011011", 18192 => "1101101011010011", 18193 => "1011001001011100", 18194 => "0011000111000111", 18195 => "1011101111000110", 18196 => "0100101111101110", 18197 => "1011011101110000", 18198 => "1110000001111011", 18199 => "0100110011111011", 18200 => "1101010101001010", 18201 => "1100011000101111", 18202 => "0101110111110011", 18203 => "0000011000001000", 18204 => "0101010111111110", 18205 => "0000001111011001", 18206 => "0111101111010110", 18207 => "1010000010001101", 18208 => "1000111111110110", 18209 => "0101000000100001", 18210 => "0011100100110010", 18211 => "1100011011011100", 18212 => "1100010101010001", 18213 => "1010100111100010", 18214 => "1101110110011011", 18215 => "0011000000110011", 18216 => "1111100101011001", 18217 => "1001000100011000", 18218 => "1111010111100111", 18219 => "0111010001011001", 18220 => "0100001111111010", 18221 => "1100011010010011", 18222 => "1010010111100010", 18223 => "1110100101011101", 18224 => "0111010101001100", 18225 => "1100000011010100", 18226 => "0011111111100110", 18227 => "1111010111011011", 18228 => "0000111110011001", 18229 => "0100100000011011", 18230 => "0011111110000100", 18231 => "1111011101010110", 18232 => "1100101001101111", 18233 => "1111110111110000", 18234 => "1100010110011001", 18235 => "0010100000111110", 18236 => "1001111000101011", 18237 => "1010101100010001", 18238 => "1000111001101010", 18239 => "1011001111011000", 18240 => "0101110100100001", 18241 => "1011011011011111", 18242 => "0111011100101111", 18243 => "0000000001101001", 18244 => "1000111110111111", 18245 => "1100111011110100", 18246 => "1100011111101110", 18247 => "1011001010110010", 18248 => "0011111001001001", 18249 => "1010101000111100", 18250 => "1111010010001111", 18251 => "0110100000000000", 18252 => "0111101101110101", 18253 => "0001110010000101", 18254 => "0101111100011010", 18255 => "0100110001111111", 18256 => "1111100110111001", 18257 => "1111000001011111", 18258 => "1110111111110111", 18259 => "0111110100111100", 18260 => "1001100001000001", 18261 => "0010010110000101", 18262 => "1001100100101110", 18263 => "1000001101101111", 18264 => "1101011101101111", 18265 => "1110000000111110", 18266 => "0010011011101101", 18267 => "0011000101000101", 18268 => "0011001101100011", 18269 => "0110010100100110", 18270 => "0001110100001100", 18271 => "1010000100010110", 18272 => "1011011101000011", 18273 => "0111001011011001", 18274 => "1000110100111100", 18275 => "0100000111110100", 18276 => "0100011111010011", 18277 => "0110110111101000", 18278 => "1101100100001011", 18279 => "1101010001001000", 18280 => "1011011101001000", 18281 => "1010001011010000", 18282 => "0011000110110100", 18283 => "0010010111110001", 18284 => "1101000011110111", 18285 => "1110111000001110", 18286 => "0010010001101000", 18287 => "0001011010001000", 18288 => "0111110001111101", 18289 => "0011001111111111", 18290 => "1010110101001100", 18291 => "1111101100100011", 18292 => "0010101010110001", 18293 => "0110111000011110", 18294 => "1000000010110000", 18295 => "1111010100010101", 18296 => "0101000110111010", 18297 => "1000101010111110", 18298 => "0100110111001100", 18299 => "0111100001010001", 18300 => "0100000101101011", 18301 => "0001110001110001", 18302 => "1111110001010111", 18303 => "0101111010001101", 18304 => "0101011001000100", 18305 => "0111010100011000", 18306 => "1110000101011010", 18307 => "0111000011010100", 18308 => "0100101010101110", 18309 => "0101010011111011", 18310 => "0001011111111111", 18311 => "0111010011111101", 18312 => "1010111101101110", 18313 => "0100100110001100", 18314 => "1001011000000011", 18315 => "0100100111100110", 18316 => "0010000011010101", 18317 => "0111101010110011", 18318 => "0010110111000011", 18319 => "1000100001010111", 18320 => "1111111101010000", 18321 => "1010010101000111", 18322 => "1011110000110001", 18323 => "1111111101100100", 18324 => "1100101111100101", 18325 => "0101011011010110", 18326 => "0000111110100011", 18327 => "1000111100011001", 18328 => "0110100011011111", 18329 => "0001001010110101", 18330 => "0011111000010010", 18331 => "0101110001010101", 18332 => "1100001011101001", 18333 => "1011011011110111", 18334 => "0111100011001000", 18335 => "0010101110010100", 18336 => "0111001001001101", 18337 => "0000110101011100", 18338 => "0101001101011110", 18339 => "1000001011001111", 18340 => "0000010000001100", 18341 => "1011011100100100", 18342 => "0011001001010110", 18343 => "1101100000010011", 18344 => "1000110111011000", 18345 => "0001100001100100", 18346 => "1110100011101001", 18347 => "0100001100001011", 18348 => "1010101100011111", 18349 => "1011110011101110", 18350 => "1110101101100010", 18351 => "1000111100110111", 18352 => "1010001010110111", 18353 => "0110000110110001", 18354 => "1001000001100100", 18355 => "0101111110001101", 18356 => "0111010011010001", 18357 => "1010110001010000", 18358 => "1111000101110010", 18359 => "1000001011010110", 18360 => "1011101101011101", 18361 => "0110011100001010", 18362 => "1001100001001001", 18363 => "1000001010111111", 18364 => "1011110000001011", 18365 => "1011000011111010", 18366 => "0000000010011010", 18367 => "0001100001011100", 18368 => "1110101010110101", 18369 => "0000000110110010", 18370 => "0010110101110001", 18371 => "0011010100010010", 18372 => "0011000011100101", 18373 => "0111010001001111", 18374 => "1000111010001000", 18375 => "1111011010000111", 18376 => "1101010011110001", 18377 => "0001101110101011", 18378 => "0111100010111011", 18379 => "1101001110101011", 18380 => "0011010010010100", 18381 => "0011111001010100", 18382 => "1111011010111111", 18383 => "0010110110110011", 18384 => "0110110011101000", 18385 => "0111010110000010", 18386 => "0001001111010100", 18387 => "0000000010010000", 18388 => "1110110011011000", 18389 => "1011100011000111", 18390 => "1100000011010101", 18391 => "0000111010011110", 18392 => "1101011000000011", 18393 => "1101000100111111", 18394 => "1000010111011110", 18395 => "1111001110001000", 18396 => "1111110110001111", 18397 => "1001011010110001", 18398 => "1000100101010101", 18399 => "1011111001010100", 18400 => "0011011011101100", 18401 => "0001011011011101", 18402 => "1110010101011111", 18403 => "0101000110110111", 18404 => "1000111100100010", 18405 => "0001110101010110", 18406 => "0011011000001100", 18407 => "1000110001111000", 18408 => "1001101110100001", 18409 => "0011001111101110", 18410 => "0010111101101110", 18411 => "1101000001111001", 18412 => "0010110011110101", 18413 => "0100001100110000", 18414 => "1111100100101100", 18415 => "0111100001001111", 18416 => "1101011010111000", 18417 => "1100100001111001", 18418 => "0010011001001111", 18419 => "1111101100010110", 18420 => "1100011000101110", 18421 => "0010011100110010", 18422 => "1101110101010001", 18423 => "1000001100110111", 18424 => "0101101110111100", 18425 => "0001010110001011", 18426 => "1000001110101001", 18427 => "0110111011110010", 18428 => "0011111101011010", 18429 => "1000000001100101", 18430 => "1101011010011110", 18431 => "1100100101001000", 18432 => "1000100010001011", 18433 => "0001011111110101", 18434 => "0000000011001010", 18435 => "1110100000011000", 18436 => "0100001011000000", 18437 => "0011011001010010", 18438 => "0100000011111110", 18439 => "0001100100101111", 18440 => "0101100000010001", 18441 => "1010000000010010", 18442 => "0001110110011111", 18443 => "0000000011111110", 18444 => "0000001011001001", 18445 => "1101100101011111", 18446 => "0011100110011101", 18447 => "1111001111010011", 18448 => "0000101011010101", 18449 => "0100110110010110", 18450 => "0000010100100011", 18451 => "1101011010111101", 18452 => "1010010000110011", 18453 => "1011011010011010", 18454 => "1110110110111000", 18455 => "0011110100110001", 18456 => "0000011110001000", 18457 => "1111100101010101", 18458 => "0101110101011100", 18459 => "1100111101110111", 18460 => "1011010010101001", 18461 => "0101011011000110", 18462 => "1011101100111011", 18463 => "1011100110110100", 18464 => "0111010110111001", 18465 => "0101011011010100", 18466 => "1111101100011111", 18467 => "1011110000100101", 18468 => "0110101110000111", 18469 => "1100111011100111", 18470 => "0011010111001010", 18471 => "0010011001001010", 18472 => "1001010010110011", 18473 => "1110001000010111", 18474 => "1110011101000000", 18475 => "1100100101010000", 18476 => "1110011000101101", 18477 => "0011100111001110", 18478 => "0101101010100110", 18479 => "0110010011001100", 18480 => "0000101011001101", 18481 => "1001110011101001", 18482 => "1101000101000111", 18483 => "0001000001001001", 18484 => "0111001101110101", 18485 => "0010011110001010", 18486 => "0101001001100100", 18487 => "0100111100000000", 18488 => "1010101000110010", 18489 => "0101011011111011", 18490 => "1011101110100101", 18491 => "1000001100111000", 18492 => "1001100000100100", 18493 => "0101101110101111", 18494 => "1000011011101101", 18495 => "1111101100010001", 18496 => "0010101010001101", 18497 => "0011011110001001", 18498 => "0011011110100010", 18499 => "0000010010111000", 18500 => "0000110111111100", 18501 => "0100110000111001", 18502 => "0101101100011011", 18503 => "1100001010101111", 18504 => "0000010110110000", 18505 => "0100101010000000", 18506 => "1111010000110100", 18507 => "0001011000101000", 18508 => "0000100010110001", 18509 => "1000111101100010", 18510 => "1010010000100001", 18511 => "0111001101000010", 18512 => "1011111101011010", 18513 => "1110011110111010", 18514 => "1010100010111001", 18515 => "0001011000100110", 18516 => "0110010000100001", 18517 => "1001100110010100", 18518 => "0110101000110101", 18519 => "1111111010110111", 18520 => "0010110111100011", 18521 => "1000111000101001", 18522 => "0101100010001101", 18523 => "0001111101111110", 18524 => "0010100100100100", 18525 => "0000100001001111", 18526 => "1111101010001010", 18527 => "1101001011100111", 18528 => "1101000100110000", 18529 => "1101101110000110", 18530 => "0110010000010111", 18531 => "1110001001000011", 18532 => "1010101011000110", 18533 => "1000101110001101", 18534 => "1010100110010001", 18535 => "0000010000010001", 18536 => "0001000011011010", 18537 => "0100000110010001", 18538 => "1011000101110011", 18539 => "0110110011000100", 18540 => "1011001101101010", 18541 => "0111110111000101", 18542 => "1110000111101110", 18543 => "1100000111110100", 18544 => "1111110110011001", 18545 => "1110111110111000", 18546 => "0110101110111100", 18547 => "1110000100110100", 18548 => "1100110010011110", 18549 => "0001001011001101", 18550 => "1001100000000010", 18551 => "0011010101011101", 18552 => "0011010110000111", 18553 => "0011100010011111", 18554 => "0001101000010010", 18555 => "0011110000111001", 18556 => "1001100111000001", 18557 => "1000000101000000", 18558 => "1000001010010111", 18559 => "0011011001010011", 18560 => "0101000011011000", 18561 => "0000010011010010", 18562 => "1101100001101101", 18563 => "1000011101001011", 18564 => "0011001110001101", 18565 => "1001110000000111", 18566 => "0110110000110011", 18567 => "1000011101000101", 18568 => "1011111010111000", 18569 => "1101111100100110", 18570 => "0010100001101110", 18571 => "1011101111011001", 18572 => "0110110011010011", 18573 => "0101111100010000", 18574 => "0000000101001010", 18575 => "0111000001100001", 18576 => "1101011111000011", 18577 => "0000111100010011", 18578 => "1000111111001010", 18579 => "1111101101011011", 18580 => "1101101011000100", 18581 => "0111100011100011", 18582 => "1111010110110010", 18583 => "0110000010110010", 18584 => "1101111011000001", 18585 => "0010110100111110", 18586 => "0000001100100001", 18587 => "0010101110010000", 18588 => "0100100111001001", 18589 => "0011010101011101", 18590 => "1101001110111000", 18591 => "0111011110010010", 18592 => "1011101110011011", 18593 => "1010011000110101", 18594 => "0011100101000101", 18595 => "0001100001100001", 18596 => "1010100011000000", 18597 => "1000001010010101", 18598 => "0011101001110101", 18599 => "1011001100110100", 18600 => "1111001100111100", 18601 => "0100001101101100", 18602 => "0010100000100000", 18603 => "0001000111111110", 18604 => "0001000000100001", 18605 => "1000010001001111", 18606 => "0100000100111011", 18607 => "1111111110011111", 18608 => "1010011110100010", 18609 => "0111100101110101", 18610 => "1101010011000100", 18611 => "0100110101010110", 18612 => "1010100110100100", 18613 => "0110101100100111", 18614 => "1010010100101111", 18615 => "0101110101001000", 18616 => "0101101000100101", 18617 => "0001100111100101", 18618 => "1011000000001101", 18619 => "1011110100101110", 18620 => "0110000010000111", 18621 => "0001100111111110", 18622 => "1000001011010000", 18623 => "1101100001100011", 18624 => "0111111000101101", 18625 => "1110011010101110", 18626 => "0010110010110000", 18627 => "0001010001010001", 18628 => "0110110001111011", 18629 => "1101011011111001", 18630 => "0001110100111111", 18631 => "1000100110000111", 18632 => "0010110000010010", 18633 => "1111000110111010", 18634 => "0001001100000001", 18635 => "1111001101101111", 18636 => "0100100111010000", 18637 => "1100001001100110", 18638 => "1011100111001101", 18639 => "1100111101011100", 18640 => "1101010011110110", 18641 => "0110111000110111", 18642 => "0101011101101010", 18643 => "0011010000101010", 18644 => "1001001111011011", 18645 => "1010101101101001", 18646 => "0110011111001000", 18647 => "1101001100110101", 18648 => "0010001000101101", 18649 => "0010000111110011", 18650 => "1100001010011110", 18651 => "1011010001110101", 18652 => "1000001011010010", 18653 => "1010100001111111", 18654 => "1000011000011011", 18655 => "0111111010100101", 18656 => "1001110001010000", 18657 => "0011010111011111", 18658 => "1000001010100011", 18659 => "1010111101011001", 18660 => "1111000101110101", 18661 => "1000110010010001", 18662 => "1011010000101001", 18663 => "1101111110101110", 18664 => "1000100111101110", 18665 => "1111001000010010", 18666 => "1100010001101001", 18667 => "1001010011110110", 18668 => "0100011000111101", 18669 => "0010000001110111", 18670 => "1001011100100000", 18671 => "1001100111111000", 18672 => "1100101000100111", 18673 => "1111110100000111", 18674 => "0010110000000100", 18675 => "0100100001110011", 18676 => "0000011100111100", 18677 => "0010011101011100", 18678 => "0001111011101110", 18679 => "0011101111001010", 18680 => "1110111101001010", 18681 => "1010110100110101", 18682 => "0100101101011111", 18683 => "1100101110100001", 18684 => "1111010101110100", 18685 => "1010101011010010", 18686 => "1001111111000101", 18687 => "1011011111010110", 18688 => "0111110001100100", 18689 => "0111011010000010", 18690 => "0000010111011100", 18691 => "0100110010001100", 18692 => "1011011010011001", 18693 => "0010110101000001", 18694 => "0000110000101010", 18695 => "1010001100101100", 18696 => "1001011111100110", 18697 => "0011011101101011", 18698 => "0101101000001011", 18699 => "0001001101111011", 18700 => "0010110100110100", 18701 => "1100001110001100", 18702 => "0001110111110000", 18703 => "1011011000101010", 18704 => "0011001101101111", 18705 => "1010010001001100", 18706 => "0101110101100010", 18707 => "1010010000101110", 18708 => "0000001110100111", 18709 => "1010001010000010", 18710 => "1101001010111000", 18711 => "0010010100001001", 18712 => "0110001001111101", 18713 => "0110100010000110", 18714 => "1010110100001011", 18715 => "0110010101101010", 18716 => "0110100001110010", 18717 => "1011111011011010", 18718 => "0000110100001000", 18719 => "0101101110101111", 18720 => "0101001111001100", 18721 => "1001000101010100", 18722 => "1110110111100011", 18723 => "1001011111010111", 18724 => "0001110101100100", 18725 => "1001011011011101", 18726 => "1011000011011110", 18727 => "0100000100101000", 18728 => "0110011101101000", 18729 => "1111010100110000", 18730 => "1100000110100110", 18731 => "1100111001010010", 18732 => "0011110111011011", 18733 => "1111010001101011", 18734 => "1101011111001011", 18735 => "1011011111101111", 18736 => "1011001010001100", 18737 => "0001100111101010", 18738 => "1100111101110001", 18739 => "0110111111000101", 18740 => "0000111110100101", 18741 => "0110001000010111", 18742 => "1000101011011110", 18743 => "1000001011010101", 18744 => "0101011101001100", 18745 => "0101010110101101", 18746 => "0010010010100110", 18747 => "0110000100011010", 18748 => "0001010100011100", 18749 => "1101001101111101", 18750 => "1001110111111100", 18751 => "1011010100001111", 18752 => "1100011101100011", 18753 => "0110011011000000", 18754 => "0010011011110000", 18755 => "1111110110100000", 18756 => "1010000111001101", 18757 => "1111001101010011", 18758 => "1011100010110100", 18759 => "0011111001101111", 18760 => "0111001100001111", 18761 => "0100110110011000", 18762 => "1110101110110100", 18763 => "0001010011110100", 18764 => "0010101010000011", 18765 => "0101111111000000", 18766 => "0010101010000101", 18767 => "0110011111101101", 18768 => "1000000000010000", 18769 => "1100001111001100", 18770 => "1010011011001101", 18771 => "0111011000001100", 18772 => "1001010010101100", 18773 => "1110111101111001", 18774 => "1010110110100001", 18775 => "1101000000110110", 18776 => "1110010010011010", 18777 => "1011000111111111", 18778 => "0100100111010110", 18779 => "0000111010001001", 18780 => "0000000111001001", 18781 => "1100010111100110", 18782 => "1100111110010110", 18783 => "0100110101100101", 18784 => "1111100000111011", 18785 => "0111010110000010", 18786 => "0010011101100010", 18787 => "1110010001101111", 18788 => "0111000111110000", 18789 => "0011010100111111", 18790 => "1010011101101001", 18791 => "0000011010100010", 18792 => "1011011010010100", 18793 => "1101010001011111", 18794 => "0100010010000000", 18795 => "1010100110110110", 18796 => "1111000010111111", 18797 => "1001110110100011", 18798 => "1111010110010111", 18799 => "1010000001101010", 18800 => "0001000011001100", 18801 => "0010111010110101", 18802 => "0011001101111011", 18803 => "1101000111001010", 18804 => "0101100000110101", 18805 => "1010101011100100", 18806 => "1111111001010100", 18807 => "1011111110100101", 18808 => "0011010101101111", 18809 => "1011110011110111", 18810 => "1111111100100000", 18811 => "1000101010110101", 18812 => "0100011011011100", 18813 => "1001110000110100", 18814 => "0110101100010001", 18815 => "0000001100001011", 18816 => "1011000011000010", 18817 => "0001010101000100", 18818 => "1110100001000001", 18819 => "1011011011101001", 18820 => "0110100111100111", 18821 => "0100110110000000", 18822 => "0001011101100011", 18823 => "0010000100111100", 18824 => "0101011001101010", 18825 => "0100010010011000", 18826 => "1101010101010100", 18827 => "1100110010010001", 18828 => "0110010101100101", 18829 => "0011110101000001", 18830 => "1000110010110101", 18831 => "1000011111101000", 18832 => "0010101111010011", 18833 => "1110101011010010", 18834 => "0001101001101011", 18835 => "0110100000111001", 18836 => "1001010111111101", 18837 => "0000000001000100", 18838 => "0011011100111011", 18839 => "0100011100011010", 18840 => "0010000000001111", 18841 => "1010010100011110", 18842 => "1011000101000001", 18843 => "1110011011111110", 18844 => "1011011100000100", 18845 => "1100011011001011", 18846 => "0101111101100001", 18847 => "1110001110011100", 18848 => "1000111101011001", 18849 => "1100010000011010", 18850 => "1111110011101110", 18851 => "0110010001100011", 18852 => "1101001011001101", 18853 => "0010011111000100", 18854 => "1110010000100110", 18855 => "0001110100010010", 18856 => "1100010010010010", 18857 => "0011111001001100", 18858 => "1000001101001101", 18859 => "0000111111101000", 18860 => "0010101100111110", 18861 => "1010101111111111", 18862 => "0110011110110010", 18863 => "0101101101111111", 18864 => "1010101110101001", 18865 => "1100011110101111", 18866 => "0011100101100100", 18867 => "1101111110001011", 18868 => "1010110001110111", 18869 => "0011100100111001", 18870 => "0011110000100001", 18871 => "1110011111001000", 18872 => "1011000101111101", 18873 => "0011100011000001", 18874 => "1010101111100011", 18875 => "0111001111000110", 18876 => "1110001000011111", 18877 => "0101000101100100", 18878 => "1011010111010011", 18879 => "1001111010000011", 18880 => "0010101100111011", 18881 => "1010000010011110", 18882 => "1000101011110000", 18883 => "1101001100000000", 18884 => "0011000010100111", 18885 => "1000110001011001", 18886 => "0100100001010011", 18887 => "0000000001001110", 18888 => "0011001011000110", 18889 => "1111011001111110", 18890 => "0000110010110010", 18891 => "0000001110111010", 18892 => "1110111001101111", 18893 => "0011100001100011", 18894 => "0110110001001000", 18895 => "1100100001101011", 18896 => "1100111001101011", 18897 => "1000011000101011", 18898 => "1010000001110010", 18899 => "0101001001010110", 18900 => "0001111111010000", 18901 => "0101011111011010", 18902 => "1110110000101011", 18903 => "1001001111101011", 18904 => "1000111111001100", 18905 => "1110111011001100", 18906 => "0000001110010101", 18907 => "1100100111101110", 18908 => "0101001101001010", 18909 => "0100111001011110", 18910 => "0010111101000001", 18911 => "1010101010101000", 18912 => "1101100010011011", 18913 => "1011100010000100", 18914 => "0011110000110011", 18915 => "0000111010111010", 18916 => "1110101011101011", 18917 => "1111011000101101", 18918 => "0111101001110111", 18919 => "0101100100101010", 18920 => "0111110000011011", 18921 => "1100011101110110", 18922 => "1010110100011011", 18923 => "1100111001010011", 18924 => "1110001001101101", 18925 => "0111001011000101", 18926 => "1010111001110010", 18927 => "1100011110110111", 18928 => "1010011101111010", 18929 => "0010010111011000", 18930 => "0111101011000110", 18931 => "0110000000111111", 18932 => "1100110111100110", 18933 => "1101110011001011", 18934 => "1101000001001001", 18935 => "1011001000111001", 18936 => "0010011010011101", 18937 => "0000100001011111", 18938 => "1100001111110110", 18939 => "1010011001011101", 18940 => "0011011111101100", 18941 => "1010000110110101", 18942 => "1010100010100011", 18943 => "0111100110000101", 18944 => "0001111001101101", 18945 => "0010001101010100", 18946 => "1100000010010011", 18947 => "1111110010000001", 18948 => "1010110001011110", 18949 => "0100111100100011", 18950 => "1111010110110100", 18951 => "1000000100011011", 18952 => "0000100011001101", 18953 => "0110000010101100", 18954 => "1010010111001011", 18955 => "0011100000110000", 18956 => "0101111101010101", 18957 => "0011010110010100", 18958 => "0110100110100010", 18959 => "1101011011100111", 18960 => "0111101101101111", 18961 => "1101100100100110", 18962 => "0110111110100110", 18963 => "0001110010110101", 18964 => "1111101011000000", 18965 => "1010101011101000", 18966 => "1110100000110000", 18967 => "1000100101111110", 18968 => "1101110100111100", 18969 => "0110001000010001", 18970 => "1111010111000001", 18971 => "1101011111100111", 18972 => "0000100110010100", 18973 => "0100000010010010", 18974 => "1011100111000110", 18975 => "0111011011101101", 18976 => "1101111011101001", 18977 => "1011011101101011", 18978 => "0110111000111010", 18979 => "0011010110101110", 18980 => "0001000110011110", 18981 => "0101110000101110", 18982 => "0000001101101010", 18983 => "1000110010010011", 18984 => "0101100101000011", 18985 => "1101001101010010", 18986 => "1000001100101000", 18987 => "1110110101110011", 18988 => "0001000011111001", 18989 => "1000010110101110", 18990 => "0000100011111010", 18991 => "1110110001100101", 18992 => "0110101011001000", 18993 => "1011010101010111", 18994 => "0010100001000011", 18995 => "0000000011000011", 18996 => "0110000110011001", 18997 => "0101100011101111", 18998 => "1110111111100100", 18999 => "1111101101100100", 19000 => "0100000110111101", 19001 => "0101110100100110", 19002 => "1010000111100000", 19003 => "1111111000010111", 19004 => "1100110010111001", 19005 => "1001101011111001", 19006 => "0011011101010010", 19007 => "1101010101010100", 19008 => "1011011110111001", 19009 => "0110111000100000", 19010 => "1111011110010111", 19011 => "1101011111000001", 19012 => "1100110001111110", 19013 => "1110111110111101", 19014 => "0111110011010010", 19015 => "1111001111101100", 19016 => "0001110100110011", 19017 => "1000101111001111", 19018 => "0101110010101010", 19019 => "1101100010001011", 19020 => "1111011000010111", 19021 => "1010101010010010", 19022 => "1000001111011000", 19023 => "0101101001111001", 19024 => "1011100010011100", 19025 => "0001100011110011", 19026 => "1111000001000000", 19027 => "0101101001110100", 19028 => "0001010100011111", 19029 => "0110001000101001", 19030 => "1010001001110010", 19031 => "0100111100011000", 19032 => "0001110011101011", 19033 => "0111000110001000", 19034 => "0010010001001110", 19035 => "1000110011101010", 19036 => "0100000101101010", 19037 => "0011010011111000", 19038 => "0010100011001000", 19039 => "1010010001011101", 19040 => "1010011010101011", 19041 => "1100011011001111", 19042 => "1011010000101100", 19043 => "1000000000111110", 19044 => "1010110100100100", 19045 => "1001001000010101", 19046 => "0010110100000110", 19047 => "0101001010010010", 19048 => "1000101000001010", 19049 => "0000000101000110", 19050 => "0100100000000110", 19051 => "0111101011010001", 19052 => "0111110010110000", 19053 => "0101010010001010", 19054 => "0111001000011110", 19055 => "0111110100010100", 19056 => "0110011110101011", 19057 => "0000000001100000", 19058 => "1101101010111000", 19059 => "1111001100000111", 19060 => "0100000101110001", 19061 => "1011111010011000", 19062 => "1000101001011111", 19063 => "1001011010100101", 19064 => "0000001111000000", 19065 => "0010100110001000", 19066 => "0101111000111011", 19067 => "0110100000111111", 19068 => "1111110011001111", 19069 => "1001110111010110", 19070 => "0001111001010110", 19071 => "1110111000110100", 19072 => "1010101000111110", 19073 => "0110000000111000", 19074 => "0000001010000001", 19075 => "1010000010110100", 19076 => "0110011010001100", 19077 => "1101110110010001", 19078 => "0010011000110001", 19079 => "1010111001111011", 19080 => "1010001101111010", 19081 => "0001001111011101", 19082 => "1110101000001101", 19083 => "1001010010111110", 19084 => "1001001010011111", 19085 => "0100101001001100", 19086 => "1101010100110111", 19087 => "0101011101001011", 19088 => "0111110110111110", 19089 => "0100001010010010", 19090 => "0001001000001101", 19091 => "1101000010010000", 19092 => "0110110010011010", 19093 => "0010001101100111", 19094 => "1101001111011001", 19095 => "0100010000100110", 19096 => "1011001000111101", 19097 => "0100100011111001", 19098 => "0101011010110100", 19099 => "0100111001101001", 19100 => "1110100111100011", 19101 => "1111000110100100", 19102 => "1010011000011110", 19103 => "1000101010001011", 19104 => "1010010111100000", 19105 => "0110001100001010", 19106 => "0000111100010000", 19107 => "1000110111011001", 19108 => "1010011001000010", 19109 => "1110100111100100", 19110 => "0001101011110011", 19111 => "1111010100000001", 19112 => "0000000000000110", 19113 => "1111010111110010", 19114 => "0010011100110001", 19115 => "1011100111100110", 19116 => "1011101101111101", 19117 => "0001100111100101", 19118 => "1111100110111100", 19119 => "1011111000101111", 19120 => "1111001000111000", 19121 => "0101101110101010", 19122 => "0000110011100111", 19123 => "0000101110100101", 19124 => "0101111010100001", 19125 => "0111110101011110", 19126 => "1100010101100001", 19127 => "1010010101111000", 19128 => "1010010100101001", 19129 => "0010100001100111", 19130 => "1111101101001101", 19131 => "1001011001110100", 19132 => "0000010110100100", 19133 => "0100101000111111", 19134 => "1100100110011000", 19135 => "1000000001111000", 19136 => "0110000011110001", 19137 => "0001000110010111", 19138 => "0000000100001111", 19139 => "0001111100111001", 19140 => "0011000000011100", 19141 => "0101000010001001", 19142 => "0011101000110111", 19143 => "1001010001010110", 19144 => "1101011101100011", 19145 => "0101100001100010", 19146 => "1111100101011001", 19147 => "1100111111011101", 19148 => "0001001000001010", 19149 => "1000001011000000", 19150 => "0101000110001001", 19151 => "1111001101100110", 19152 => "1101110011100100", 19153 => "1000101011100100", 19154 => "0111001111011010", 19155 => "0110110010010010", 19156 => "0110111111000000", 19157 => "0001110111111010", 19158 => "0111001001011010", 19159 => "1101010001110001", 19160 => "1010001010011001", 19161 => "0001110000110110", 19162 => "1111111010001101", 19163 => "1001011101000110", 19164 => "0010001110001011", 19165 => "0000101011001110", 19166 => "1110110101100010", 19167 => "1011001111011011", 19168 => "0100001100000001", 19169 => "0111110100110011", 19170 => "1011101110000110", 19171 => "1100111000011001", 19172 => "1100110010110101", 19173 => "0101011111110110", 19174 => "1111111100101101", 19175 => "0101110100000010", 19176 => "0000001111000110", 19177 => "0101100001101000", 19178 => "1111111111111110", 19179 => "1110101011001000", 19180 => "0101001101001101", 19181 => "0101001110001011", 19182 => "1100000101010010", 19183 => "1001111011110011", 19184 => "1011111000111100", 19185 => "1000101100101100", 19186 => "0100010001111000", 19187 => "1000000111100110", 19188 => "0101111000011001", 19189 => "1100000111101011", 19190 => "1111000011000100", 19191 => "1010111111110111", 19192 => "1000110001110111", 19193 => "1111011101011011", 19194 => "0110010000011011", 19195 => "0110101101001000", 19196 => "0010001111101010", 19197 => "1011000110100101", 19198 => "1110011010110001", 19199 => "0000110001001011", 19200 => "0110010111101110", 19201 => "0110110001100010", 19202 => "0110011001011011", 19203 => "0011110110000000", 19204 => "1111111110101011", 19205 => "0011000101000010", 19206 => "0111011000101001", 19207 => "1110001100011011", 19208 => "1101101110001100", 19209 => "0111010001001010", 19210 => "0001001100011101", 19211 => "0010001001101101", 19212 => "0010011100101010", 19213 => "1101101111101110", 19214 => "1110001001100111", 19215 => "1001110011110110", 19216 => "0011010101011001", 19217 => "0011001111001111", 19218 => "0000000010001101", 19219 => "1011010101110101", 19220 => "1101101110101000", 19221 => "1100010110111100", 19222 => "1010101001000001", 19223 => "1110011101000010", 19224 => "0010010001010001", 19225 => "0010010110010010", 19226 => "1110101000011010", 19227 => "1010111010111111", 19228 => "0011011110010111", 19229 => "1110001110010011", 19230 => "1010001110110000", 19231 => "0010000100110111", 19232 => "1111000000101010", 19233 => "0101001101100110", 19234 => "0011000000111000", 19235 => "1000111001110101", 19236 => "1010101101101001", 19237 => "1010101000100000", 19238 => "0101000011100100", 19239 => "1000000101011011", 19240 => "0001001000101110", 19241 => "0111001010100111", 19242 => "1010011011110111", 19243 => "0110110111110010", 19244 => "0001010011101101", 19245 => "1101110110111011", 19246 => "1101000111101111", 19247 => "1101100011000111", 19248 => "1100000111100001", 19249 => "0100110100010010", 19250 => "0011100100110010", 19251 => "1110000110000010", 19252 => "0010100100111110", 19253 => "1111001001101011", 19254 => "0000010111100000", 19255 => "1101000100100110", 19256 => "1101100011110000", 19257 => "0110010111010111", 19258 => "0100100101111110", 19259 => "1100000001111111", 19260 => "1000100001110001", 19261 => "1011011100011001", 19262 => "0101011010010010", 19263 => "0000001111101100", 19264 => "0000111110001111", 19265 => "1100110000010101", 19266 => "1100101000101101", 19267 => "0101111111000000", 19268 => "0001000001000111", 19269 => "1110011011100010", 19270 => "1100100111100010", 19271 => "1010100010001010", 19272 => "0001100011011111", 19273 => "0001111000011001", 19274 => "1100010010100010", 19275 => "1011010011111110", 19276 => "1001001111011100", 19277 => "1100110111110011", 19278 => "0011110001001101", 19279 => "1101101000010101", 19280 => "1010100101110010", 19281 => "0110110101101100", 19282 => "0110111100001100", 19283 => "1000101001110100", 19284 => "1000110011000110", 19285 => "0000110001000110", 19286 => "1100001000010011", 19287 => "0011100010100000", 19288 => "0010011110000111", 19289 => "0001110110011001", 19290 => "0000110100000111", 19291 => "1101000111000010", 19292 => "1010000101001001", 19293 => "1110101010101000", 19294 => "0000001110101101", 19295 => "0011011100000011", 19296 => "1100000100111101", 19297 => "1001000111110110", 19298 => "0101100101100011", 19299 => "0000100001000001", 19300 => "0000111000001011", 19301 => "1011010011100100", 19302 => "0000000101011000", 19303 => "0011000000110110", 19304 => "0001001111011011", 19305 => "1111000001110111", 19306 => "1101111101110100", 19307 => "1010101011101010", 19308 => "0100000100111000", 19309 => "0010111101001100", 19310 => "1110110111011100", 19311 => "0111110101000001", 19312 => "1001110111111011", 19313 => "1011100110010010", 19314 => "0011100101100101", 19315 => "0000001001000101", 19316 => "0010100000010011", 19317 => "0000110111001001", 19318 => "1101000111101100", 19319 => "0101110101110100", 19320 => "1101110011101001", 19321 => "0000000010111101", 19322 => "1100101010101001", 19323 => "1010010001111100", 19324 => "0110001111001000", 19325 => "0100111110010111", 19326 => "0010010010011100", 19327 => "0000000010110011", 19328 => "0010110100111110", 19329 => "1101111010000001", 19330 => "1101011001110000", 19331 => "0010011110100010", 19332 => "1110010100010001", 19333 => "0011011001111111", 19334 => "1111010000110000", 19335 => "0110110101101010", 19336 => "1110111110001111", 19337 => "0001101100101110", 19338 => "0001000101110100", 19339 => "1111101110111100", 19340 => "0101011100110001", 19341 => "0011100111111000", 19342 => "0111101101000010", 19343 => "0111110000001110", 19344 => "0010100111011111", 19345 => "1101010010000010", 19346 => "0100111001010011", 19347 => "1010111110111011", 19348 => "1100110110011000", 19349 => "1001001101000101", 19350 => "1010111011101001", 19351 => "0001111100111000", 19352 => "0101110100011100", 19353 => "1100100110011011", 19354 => "0100010110100000", 19355 => "0101111101000001", 19356 => "0001011000101001", 19357 => "0100101111100100", 19358 => "0110111100000010", 19359 => "1110101010000101", 19360 => "1001011101110001", 19361 => "0001001010100110", 19362 => "1000010101010000", 19363 => "1101111000101000", 19364 => "0100010000101100", 19365 => "1001111101001000", 19366 => "0001100111000010", 19367 => "1000000010011001", 19368 => "0001001000010110", 19369 => "1100001001010010", 19370 => "0010111100011001", 19371 => "1010110101111101", 19372 => "0000000011000011", 19373 => "1001001011111010", 19374 => "0010111111011000", 19375 => "1100001001111011", 19376 => "0000011010010101", 19377 => "0100110001001110", 19378 => "1011100110111101", 19379 => "0010011101011100", 19380 => "0001101000011101", 19381 => "0001000001000110", 19382 => "1011010000110011", 19383 => "0010101111111110", 19384 => "0001100111011001", 19385 => "1100000110001111", 19386 => "1001101011011110", 19387 => "0000000100001111", 19388 => "0001000100101000", 19389 => "1010011011101010", 19390 => "1111111111101001", 19391 => "0001100111000001", 19392 => "1010110001101110", 19393 => "0001000110101111", 19394 => "1110110010010110", 19395 => "1011111011111010", 19396 => "0101111111110100", 19397 => "0001001000001111", 19398 => "0000011001101100", 19399 => "1111111110010011", 19400 => "1010110011001011", 19401 => "0101001110011111", 19402 => "0000001011101000", 19403 => "1100100101010101", 19404 => "1111111001010101", 19405 => "0011001101101010", 19406 => "0111000101111111", 19407 => "0111000010000111", 19408 => "0110000101100101", 19409 => "1010100101011100", 19410 => "1000111011111001", 19411 => "0111111110000101", 19412 => "0011101110001101", 19413 => "0011101101111011", 19414 => "1001111001101010", 19415 => "0100000011110010", 19416 => "0001011100000010", 19417 => "0000011101110110", 19418 => "0000101111010011", 19419 => "0000000101100001", 19420 => "0100110100111110", 19421 => "0110110111011100", 19422 => "0010111001100100", 19423 => "1101101001111110", 19424 => "0000110111110011", 19425 => "0010111111011111", 19426 => "0001011110000100", 19427 => "0011000001010110", 19428 => "1100010111110100", 19429 => "0110000011101101", 19430 => "0110000101010111", 19431 => "1010001010101010", 19432 => "1111111000001011", 19433 => "0000110111110101", 19434 => "0111011110110111", 19435 => "0100011001100101", 19436 => "1011010110001000", 19437 => "1000101100110010", 19438 => "1101101111111010", 19439 => "1110110100100001", 19440 => "0010001101110001", 19441 => "0101111110100100", 19442 => "1111001101010101", 19443 => "0010100000101111", 19444 => "1000101000001010", 19445 => "1001100001110000", 19446 => "1011011001101101", 19447 => "0000110101000110", 19448 => "0010010000001100", 19449 => "1100011001110111", 19450 => "0001101001011110", 19451 => "1110000110100001", 19452 => "1110010100010011", 19453 => "0111101110000101", 19454 => "0011011000110000", 19455 => "0100110100011101", 19456 => "0110111110001011", 19457 => "0101100111011010", 19458 => "0001001001110111", 19459 => "0111011101111111", 19460 => "0010011100110110", 19461 => "0000001110010010", 19462 => "0101001101111100", 19463 => "1111010011011111", 19464 => "1111000111001100", 19465 => "0111011001011011", 19466 => "1001011100101111", 19467 => "0101000101110100", 19468 => "0010011011000110", 19469 => "1011100010010000", 19470 => "1011111110110101", 19471 => "1100011111101110", 19472 => "0110100000100000", 19473 => "0011011101010110", 19474 => "1101011000111000", 19475 => "0100010111001010", 19476 => "1011001001101110", 19477 => "0101100000000000", 19478 => "0101111100101110", 19479 => "1010100101000000", 19480 => "0011100110111001", 19481 => "0011110111110110", 19482 => "0110101100111100", 19483 => "1111011011100010", 19484 => "1001101100000011", 19485 => "0000001101011100", 19486 => "0111101000000101", 19487 => "1111110001010111", 19488 => "0001111010111000", 19489 => "1101101111001010", 19490 => "0000000000001100", 19491 => "1010101100010001", 19492 => "1001010100100001", 19493 => "0111011010111011", 19494 => "1110010000010111", 19495 => "0101110010101011", 19496 => "1010000111010001", 19497 => "0100100101111110", 19498 => "1110110111111111", 19499 => "1000100001101000", 19500 => "1001110010001101", 19501 => "0001011001011101", 19502 => "0011100100000100", 19503 => "0000000000010011", 19504 => "0000010000010111", 19505 => "0110010100000101", 19506 => "0110110010110110", 19507 => "0010110110111101", 19508 => "1101011111001011", 19509 => "1111011111011111", 19510 => "1010110011010010", 19511 => "0000010110001001", 19512 => "0111111111001101", 19513 => "1101100100000001", 19514 => "1101111011010110", 19515 => "0011110101100001", 19516 => "0011100001001110", 19517 => "1010110100100101", 19518 => "0101100110001010", 19519 => "0000001101101001", 19520 => "0110011000101001", 19521 => "0110100001111100", 19522 => "1111011101011011", 19523 => "0101111000001010", 19524 => "0101000011110011", 19525 => "1010110100001001", 19526 => "0111111011001001", 19527 => "1011100000011000", 19528 => "0000011010101000", 19529 => "0111110000101110", 19530 => "1010011110101000", 19531 => "1000011011100000", 19532 => "1000000001000101", 19533 => "0101110010001111", 19534 => "1000110000100001", 19535 => "1101111111110000", 19536 => "1110011110010110", 19537 => "1101111101001010", 19538 => "0011011001001000", 19539 => "1111000101000000", 19540 => "0110010010010000", 19541 => "1101000110111001", 19542 => "0111111011010000", 19543 => "1101110010001011", 19544 => "0110101100011011", 19545 => "0010110001100011", 19546 => "0111111000110010", 19547 => "1011000111101111", 19548 => "1111110001000011", 19549 => "1100011010101001", 19550 => "0101011111011111", 19551 => "1101100010000110", 19552 => "0011100001111010", 19553 => "1100011110011000", 19554 => "0101011101101110", 19555 => "0100100100001101", 19556 => "1110010001001111", 19557 => "0010110000110010", 19558 => "0101001001110010", 19559 => "0110110011101101", 19560 => "1100011111100111", 19561 => "1010110111001100", 19562 => "1000010101000011", 19563 => "1001110010101100", 19564 => "1001111110000001", 19565 => "0011011110010111", 19566 => "0010010010110010", 19567 => "0000011111110110", 19568 => "0101011111001110", 19569 => "1000000101001000", 19570 => "0000001101100001", 19571 => "0000100101110001", 19572 => "0000110010001000", 19573 => "0010111101101101", 19574 => "0001001000000100", 19575 => "1010001110101011", 19576 => "1111000101000101", 19577 => "0011101000100110", 19578 => "1101101110001110", 19579 => "0101111110110111", 19580 => "0111001100110111", 19581 => "1110001001111111", 19582 => "1100110001000111", 19583 => "1100100101000001", 19584 => "1000001001010011", 19585 => "0100101111101101", 19586 => "1010000110100100", 19587 => "1100101011100100", 19588 => "0011001010000001", 19589 => "1011001110001110", 19590 => "1000000101011101", 19591 => "1011001001101101", 19592 => "0000011111101011", 19593 => "1100000000111111", 19594 => "0010100001111000", 19595 => "1100110100101100", 19596 => "1100010001001001", 19597 => "1111010101011100", 19598 => "1110010001101100", 19599 => "1011010101000100", 19600 => "0110101010000001", 19601 => "0111000100111100", 19602 => "1100011101000011", 19603 => "1110010000110011", 19604 => "0101100110011000", 19605 => "0011000110100111", 19606 => "0010111111101010", 19607 => "0001001001100010", 19608 => "0110100110111000", 19609 => "1101011001001100", 19610 => "1001011001001100", 19611 => "0010010001000111", 19612 => "1000111100000000", 19613 => "1110000000101001", 19614 => "0000110110110101", 19615 => "1100100001010001", 19616 => "0100111111111101", 19617 => "1001010111100010", 19618 => "0000000001101001", 19619 => "1110100100101100", 19620 => "1100011111001000", 19621 => "1001001011111100", 19622 => "0011101101000110", 19623 => "1111001001000111", 19624 => "0110111100001010", 19625 => "1110000011111000", 19626 => "1101011110100111", 19627 => "0001111010011110", 19628 => "1010000010111101", 19629 => "1100111111011110", 19630 => "1000110001000101", 19631 => "0100110001010111", 19632 => "0110111110001101", 19633 => "0001111110010011", 19634 => "1001101011101010", 19635 => "0111101011101000", 19636 => "0000101010001101", 19637 => "0110110101110000", 19638 => "1000010101000101", 19639 => "1001111010101111", 19640 => "1101000000110110", 19641 => "0101110100011100", 19642 => "1001000101000000", 19643 => "0110110110010000", 19644 => "0000001000101101", 19645 => "0111100001001000", 19646 => "0011100100111101", 19647 => "1101001100011000", 19648 => "0010011001100101", 19649 => "1001001100100010", 19650 => "1011110101001011", 19651 => "0010101000110000", 19652 => "1101011101010110", 19653 => "0110100100010001", 19654 => "0111001011111111", 19655 => "0011011101001001", 19656 => "0101110001100100", 19657 => "0110001110011111", 19658 => "0010011100001100", 19659 => "1001100010110011", 19660 => "1100010100100111", 19661 => "1101011001010101", 19662 => "0101010110001101", 19663 => "1001001101110100", 19664 => "0010111111001111", 19665 => "0011000000000100", 19666 => "1101000010010101", 19667 => "1101011111011110", 19668 => "0101011000001110", 19669 => "1010000011100011", 19670 => "1101111100000001", 19671 => "1001010100110101", 19672 => "1111010000100111", 19673 => "1111010111111011", 19674 => "0111110000110101", 19675 => "0110100001000101", 19676 => "0000000000000111", 19677 => "1111100110010101", 19678 => "0101100000111000", 19679 => "1111100000110010", 19680 => "1011100001000000", 19681 => "0100010110101110", 19682 => "0101110100100111", 19683 => "1001100000110111", 19684 => "1110001111010000", 19685 => "1100010101111101", 19686 => "1011010110011110", 19687 => "1111101011011110", 19688 => "1100111011001101", 19689 => "1110001101101001", 19690 => "0011010011110001", 19691 => "0001110110000011", 19692 => "0000110110101101", 19693 => "1010100000011010", 19694 => "1001010010101110", 19695 => "0000100010001111", 19696 => "0100110000111011", 19697 => "0100101100001110", 19698 => "0101001111110011", 19699 => "1001100010111000", 19700 => "1001100101010110", 19701 => "0101000110110110", 19702 => "0000011011011110", 19703 => "0011110101101110", 19704 => "0010100100101101", 19705 => "1100011101010110", 19706 => "1110111100110000", 19707 => "0001100111010010", 19708 => "0100010010110101", 19709 => "0011110100111011", 19710 => "1011110110010100", 19711 => "1100000110110011", 19712 => "0010001010011101", 19713 => "0110000110101100", 19714 => "1111111110001000", 19715 => "1000111010101011", 19716 => "1001000111111111", 19717 => "1000110000010100", 19718 => "0110111100111111", 19719 => "1101011101111011", 19720 => "0011000111001110", 19721 => "1011111101100011", 19722 => "1010111111011010", 19723 => "0010000010010100", 19724 => "1101101010010110", 19725 => "0010110111100010", 19726 => "1000110110011000", 19727 => "0001010010111011", 19728 => "1111100110001000", 19729 => "0011001010110101", 19730 => "1101001101110001", 19731 => "0011001111011001", 19732 => "0100001100111011", 19733 => "1110111000000001", 19734 => "0111000001001111", 19735 => "1010101010000101", 19736 => "0000011101101001", 19737 => "1111110011110101", 19738 => "0110100101111010", 19739 => "1011111111101101", 19740 => "1110110111000000", 19741 => "1100011100000010", 19742 => "0001010011101101", 19743 => "1010011110001100", 19744 => "0101000111001001", 19745 => "0001010011011000", 19746 => "1001001001111110", 19747 => "1011111101101111", 19748 => "0111001111011010", 19749 => "0010001000010010", 19750 => "0000101110111001", 19751 => "0000011011111010", 19752 => "1101101001101001", 19753 => "1100000000111001", 19754 => "1111101010100100", 19755 => "0101111001000001", 19756 => "1001110100000110", 19757 => "1011011000011110", 19758 => "0111010000000010", 19759 => "0101001010111100", 19760 => "0011010011110101", 19761 => "1001110000100100", 19762 => "0100011100011111", 19763 => "1100011010100001", 19764 => "1001111111101000", 19765 => "0111001011000000", 19766 => "1111101100010101", 19767 => "1100101100001110", 19768 => "0010010001111100", 19769 => "1011111001001001", 19770 => "1110000001110000", 19771 => "1111100010001111", 19772 => "0010010100100111", 19773 => "0111000111011110", 19774 => "0110001001110111", 19775 => "0100110101010110", 19776 => "1010000111111011", 19777 => "0001000011010000", 19778 => "0001010011011101", 19779 => "1010001110110110", 19780 => "1110110001111011", 19781 => "0111101100000010", 19782 => "1011110111001110", 19783 => "0011101100000011", 19784 => "0110111111111001", 19785 => "0000110110110010", 19786 => "0110110001010000", 19787 => "0001000110000111", 19788 => "0010001101101001", 19789 => "1110111110100101", 19790 => "1101010111000001", 19791 => "1011011101100101", 19792 => "0111001011110010", 19793 => "1011101110011111", 19794 => "1100000111111111", 19795 => "1001010101110101", 19796 => "1110001110001110", 19797 => "0110001001010110", 19798 => "1101100111011010", 19799 => "0101011100111011", 19800 => "1001000110101110", 19801 => "0100101100010000", 19802 => "0111011100011000", 19803 => "1100100001111110", 19804 => "0110011110010110", 19805 => "0100000011000101", 19806 => "0000011010100110", 19807 => "1111010000101100", 19808 => "0110000100110111", 19809 => "0011100000010010", 19810 => "1001111011011011", 19811 => "1001101011000110", 19812 => "0011110111111001", 19813 => "0101000011100111", 19814 => "1101001010010011", 19815 => "0000111001001100", 19816 => "0101100001100111", 19817 => "0110000111100001", 19818 => "1111000111110101", 19819 => "1001001010011011", 19820 => "1110100000000000", 19821 => "0101010010100101", 19822 => "1111111000001100", 19823 => "1111110111110101", 19824 => "1110111101110101", 19825 => "1011000011010000", 19826 => "0100100001100010", 19827 => "0110111000101011", 19828 => "0011100111011100", 19829 => "1101010110011111", 19830 => "0001110001001010", 19831 => "0110101111001101", 19832 => "1101100100010010", 19833 => "1110101101100101", 19834 => "0000101100101010", 19835 => "0101010011010100", 19836 => "0111000011001000", 19837 => "1001000101100111", 19838 => "1011001111110101", 19839 => "0000000100110000", 19840 => "1100000111010000", 19841 => "0111110010100011", 19842 => "1010001111100000", 19843 => "1111001000100011", 19844 => "0100100010000100", 19845 => "0100000110000110", 19846 => "1101010101110010", 19847 => "0010000001001111", 19848 => "0001000011100111", 19849 => "0101110011100001", 19850 => "0111011101110100", 19851 => "0010101100111000", 19852 => "1000010100000001", 19853 => "0100011100111110", 19854 => "0110111111100110", 19855 => "1101101101010101", 19856 => "1011010110011100", 19857 => "0100000101001111", 19858 => "0000010101111001", 19859 => "0101010001100110", 19860 => "0011101000110100", 19861 => "0100010111110111", 19862 => "0000000101000110", 19863 => "0101110111111010", 19864 => "0111101001110001", 19865 => "1110100000100011", 19866 => "0001111101100110", 19867 => "0000010110101101", 19868 => "1100101000010111", 19869 => "1100100101001011", 19870 => "0110000111100101", 19871 => "1010100111011000", 19872 => "1110000111011110", 19873 => "1000001101001010", 19874 => "1101000110100111", 19875 => "0110111100001111", 19876 => "1001000000110011", 19877 => "0010101010011010", 19878 => "1011001000001011", 19879 => "1101010101111001", 19880 => "0000010010000000", 19881 => "0001110101000011", 19882 => "0010111010010001", 19883 => "1100101101000011", 19884 => "1001111101010111", 19885 => "0011100010111001", 19886 => "1000011110000011", 19887 => "1101100010101011", 19888 => "1001101011111011", 19889 => "1011110011111011", 19890 => "0010101110100100", 19891 => "1110110101010111", 19892 => "1100010010111000", 19893 => "0000001000001010", 19894 => "0111001011101100", 19895 => "0110100001111010", 19896 => "1000000001010000", 19897 => "1011101111101101", 19898 => "0001101010100001", 19899 => "1101011111001000", 19900 => "0111110011001001", 19901 => "0001010010000110", 19902 => "0100111001101000", 19903 => "1000111010111101", 19904 => "1110111011010100", 19905 => "0110111111111011", 19906 => "1100100111111111", 19907 => "1000000011001100", 19908 => "0101100010010100", 19909 => "1100111100001010", 19910 => "1101011110000000", 19911 => "0100000011001111", 19912 => "1010100010111101", 19913 => "0110001000010111", 19914 => "1000001000011010", 19915 => "1111100110001101", 19916 => "1101101100100101", 19917 => "0110000001110010", 19918 => "0001110011100111", 19919 => "1111110111000000", 19920 => "1011010101001110", 19921 => "0010111011101111", 19922 => "0100000000110100", 19923 => "1010110010111111", 19924 => "0010001110111000", 19925 => "1010010100101010", 19926 => "0111010110111101", 19927 => "0000001011001011", 19928 => "0011110000100010", 19929 => "1001011110101011", 19930 => "0101111111011000", 19931 => "1010111101010100", 19932 => "0101101111010001", 19933 => "1001100010011111", 19934 => "1001110101000100", 19935 => "0001100111001001", 19936 => "0000010110101100", 19937 => "0011101011111101", 19938 => "1011100011100000", 19939 => "1001001100011010", 19940 => "1010010110000011", 19941 => "0111111011011110", 19942 => "1101110100010011", 19943 => "1101001110101000", 19944 => "1100001010111001", 19945 => "1001110100111011", 19946 => "1011010000100010", 19947 => "1101101101101101", 19948 => "1010110011101110", 19949 => "1110011101000011", 19950 => "0011010001111110", 19951 => "0101001110000110", 19952 => "0110010100000000", 19953 => "1000011010000110", 19954 => "1010111111100011", 19955 => "1000000010111110", 19956 => "0000010110101001", 19957 => "1100000011011000", 19958 => "0101011101100000", 19959 => "1010110100001101", 19960 => "1110101010110110", 19961 => "1010001110000101", 19962 => "1100111101010110", 19963 => "0111110100110101", 19964 => "1000100010010110", 19965 => "0110111101010100", 19966 => "0001001001010101", 19967 => "1011111100011110", 19968 => "1011101100100010", 19969 => "0000001101101100", 19970 => "0101111101101000", 19971 => "1000111001100001", 19972 => "0011100011000010", 19973 => "1000011011010101", 19974 => "0111100011101110", 19975 => "0010111111101000", 19976 => "0001011110001110", 19977 => "0010000010100001", 19978 => "1010111000100110", 19979 => "1000110101000000", 19980 => "1000100101000011", 19981 => "0001001110010010", 19982 => "1010100110110001", 19983 => "1011101111111000", 19984 => "0000011100011010", 19985 => "1110010100000001", 19986 => "0001001010111110", 19987 => "1000010110101010", 19988 => "1000111011110111", 19989 => "0100101011001000", 19990 => "0010001001011100", 19991 => "0100110011001011", 19992 => "1101001011010110", 19993 => "0011100101101001", 19994 => "1011110110111110", 19995 => "0001000011110011", 19996 => "0100100101111110", 19997 => "1001000101000001", 19998 => "0111000000000111", 19999 => "1111010010100111", 20000 => "0010001100111111", 20001 => "0101000000001010", 20002 => "0010111010100011", 20003 => "0000011001000010", 20004 => "1100000001001001", 20005 => "1011011000001101", 20006 => "0110100011010000", 20007 => "1000111000111000", 20008 => "1001001011101100", 20009 => "0010110001111100", 20010 => "0000000010011111", 20011 => "0111111000000111", 20012 => "0010100111001101", 20013 => "1011110011100111", 20014 => "0101000100100011", 20015 => "0011001101100000", 20016 => "0010111111011111", 20017 => "0010011011100110", 20018 => "1111111111011001", 20019 => "1100101011110100", 20020 => "0100101000101111", 20021 => "1000001110110101", 20022 => "1000001000110001", 20023 => "0100011011101011", 20024 => "0010010000110100", 20025 => "0101001010101111", 20026 => "0011110111101001", 20027 => "1101101011101000", 20028 => "0110001111100001", 20029 => "0011010110010101", 20030 => "0111000010110110", 20031 => "1010100001110111", 20032 => "0101011100111111", 20033 => "1110011110111001", 20034 => "0110100101001110", 20035 => "1001010010100011", 20036 => "1000111110111110", 20037 => "0111011111011101", 20038 => "1100001001101011", 20039 => "0000000111101110", 20040 => "1011000101010111", 20041 => "1001101111010001", 20042 => "0101010000001000", 20043 => "0111010101101011", 20044 => "1101000100100100", 20045 => "1011010000111001", 20046 => "1101101001000100", 20047 => "1101000110001101", 20048 => "1101111101111011", 20049 => "1110010101110000", 20050 => "0110011010000000", 20051 => "0011111101101111", 20052 => "0011111101111010", 20053 => "0011001001101111", 20054 => "0111011110011001", 20055 => "0110001110010111", 20056 => "0001100010101001", 20057 => "0110001001110111", 20058 => "0110011011111001", 20059 => "0101011000001011", 20060 => "0111110001000010", 20061 => "1101111010101100", 20062 => "0001101110101010", 20063 => "0010101000110111", 20064 => "1101010111000100", 20065 => "0111010101001000", 20066 => "0011111010110110", 20067 => "0110110100000100", 20068 => "1101001010001000", 20069 => "1100010011101100", 20070 => "1101111011001000", 20071 => "1101111110001111", 20072 => "1100001000111000", 20073 => "0100000101000110", 20074 => "1111101101000110", 20075 => "1100001000111000", 20076 => "0100100111001001", 20077 => "1001001011111000", 20078 => "1111100000101011", 20079 => "0010011101010010", 20080 => "1011111010010110", 20081 => "0100001110111001", 20082 => "0100111101110110", 20083 => "0111010101010111", 20084 => "0111110001111011", 20085 => "1001011010111001", 20086 => "0111110110010110", 20087 => "0001000111010110", 20088 => "0001100000110101", 20089 => "1100111100011000", 20090 => "1000100001110110", 20091 => "0110010100100011", 20092 => "0111011100111011", 20093 => "0001100110000100", 20094 => "1010101000110110", 20095 => "0111011100110000", 20096 => "0101001100110111", 20097 => "1011101011001110", 20098 => "1111101110001110", 20099 => "1010101001010010", 20100 => "1101001011010111", 20101 => "1100101111100010", 20102 => "1001110001010111", 20103 => "1001000100000010", 20104 => "1010011001110111", 20105 => "1110011111000010", 20106 => "1001111010000101", 20107 => "1000101011111110", 20108 => "1010010100000100", 20109 => "1101101011011110", 20110 => "0100000101111110", 20111 => "1001001111100110", 20112 => "1010010011100000", 20113 => "0010110011000100", 20114 => "1001100110011010", 20115 => "0000001010110100", 20116 => "1000010100100110", 20117 => "0100010010011011", 20118 => "0000101001111110", 20119 => "0010000000001001", 20120 => "1111111001001001", 20121 => "0110101111010010", 20122 => "0001111001110011", 20123 => "1111001110000011", 20124 => "1110111111101101", 20125 => "1010110001111010", 20126 => "0111011011111010", 20127 => "0100101011110000", 20128 => "1001101010110011", 20129 => "1011111111111101", 20130 => "0100110010011110", 20131 => "1110011111110000", 20132 => "1001110101111010", 20133 => "1101011011001010", 20134 => "1110011100100100", 20135 => "0111101011101010", 20136 => "1010000011111100", 20137 => "0101000111011100", 20138 => "1100011110111000", 20139 => "1111110001110100", 20140 => "0101111000001001", 20141 => "1001110010001001", 20142 => "1100100101011000", 20143 => "1110010101111001", 20144 => "1000001110010010", 20145 => "1000000101010110", 20146 => "1100011100111100", 20147 => "1010011010010100", 20148 => "0101110100100001", 20149 => "0011110101111101", 20150 => "1100100010101000", 20151 => "0101110101000000", 20152 => "0001101111001000", 20153 => "1011000000001101", 20154 => "0101100101100001", 20155 => "0000011111000100", 20156 => "0101010001111111", 20157 => "0111100101111101", 20158 => "1001100000000011", 20159 => "1010101010010000", 20160 => "0010011010100011", 20161 => "0111110000011101", 20162 => "0110001010111110", 20163 => "0011101001111100", 20164 => "0110111110110101", 20165 => "1010101010010111", 20166 => "1010011110110011", 20167 => "0001110111011001", 20168 => "1110001000110111", 20169 => "0011000000001000", 20170 => "1011111110001001", 20171 => "1110111000100000", 20172 => "0001001010001011", 20173 => "1100010000101011", 20174 => "0101000100011011", 20175 => "0011101100111010", 20176 => "0001111101010011", 20177 => "0110010011011101", 20178 => "0010001011010000", 20179 => "0101001011001101", 20180 => "1000010001000001", 20181 => "1111100110000011", 20182 => "0111010100010111", 20183 => "1111001110111101", 20184 => "0111110101100100", 20185 => "0100011110101110", 20186 => "0110101101000100", 20187 => "1111001110101100", 20188 => "1011011000101010", 20189 => "1111001111001010", 20190 => "1001111110110100", 20191 => "1100101010111110", 20192 => "0001001000010110", 20193 => "1001101001100010", 20194 => "1011100100001100", 20195 => "0010001101011111", 20196 => "0011000001111010", 20197 => "1001011000110101", 20198 => "0110000100110010", 20199 => "0010010111011111", 20200 => "0011000111001111", 20201 => "0000111010010000", 20202 => "0000011111010110", 20203 => "0100111010010110", 20204 => "0010011110110110", 20205 => "1100101010100011", 20206 => "0011001000101011", 20207 => "0010000001111110", 20208 => "1111011101010111", 20209 => "0000110000110001", 20210 => "0110000000110000", 20211 => "0010101000110000", 20212 => "1100001101111010", 20213 => "1110010011111001", 20214 => "1111011111010111", 20215 => "1010010111100111", 20216 => "0111011011101000", 20217 => "1111010001000011", 20218 => "0010101100101001", 20219 => "0101010000011001", 20220 => "0000001111001000", 20221 => "1000111010101101", 20222 => "0101110111111100", 20223 => "0100010000110010", 20224 => "1100001000101000", 20225 => "0100110010011011", 20226 => "1110001010110110", 20227 => "0101001100100101", 20228 => "0000101011001011", 20229 => "1000101010001101", 20230 => "1100101000001100", 20231 => "0001101111001101", 20232 => "0110111010010000", 20233 => "1100010100111100", 20234 => "1101100110101101", 20235 => "0100010001011111", 20236 => "0100000110101011", 20237 => "1100100100100100", 20238 => "1100111001000101", 20239 => "0010101100010011", 20240 => "0001010010101110", 20241 => "0110101110010110", 20242 => "1000100110010110", 20243 => "0100100011100000", 20244 => "1000100110001010", 20245 => "1010000110011101", 20246 => "0100111010011010", 20247 => "1101010110111101", 20248 => "1101010000111011", 20249 => "0000011111101111", 20250 => "1101110010000101", 20251 => "0111011011010010", 20252 => "1111110011010110", 20253 => "1110001101001000", 20254 => "1000001111101010", 20255 => "1001101010010101", 20256 => "0000111000001101", 20257 => "1001111101000001", 20258 => "0001101100111101", 20259 => "0000100000101010", 20260 => "0110100011001110", 20261 => "1110101101001000", 20262 => "1100111111100011", 20263 => "1000010101001000", 20264 => "0111000000011011", 20265 => "0110000010010011", 20266 => "1011100000100100", 20267 => "1101000111101101", 20268 => "1010100010111001", 20269 => "1001000000000010", 20270 => "0110110011101011", 20271 => "0110010010010011", 20272 => "1101010111111110", 20273 => "1110010111100000", 20274 => "1101010001111110", 20275 => "0101100110000001", 20276 => "1101000011111011", 20277 => "0100100001100100", 20278 => "0100010110010101", 20279 => "0101111001000011", 20280 => "0000000100001101", 20281 => "1101110101011000", 20282 => "0101010110101101", 20283 => "1010101011001000", 20284 => "1010000110111101", 20285 => "0111101101111010", 20286 => "0111101111011011", 20287 => "1001110001011111", 20288 => "0101101101110100", 20289 => "1001101011101001", 20290 => "0110111001001111", 20291 => "0010010010011100", 20292 => "1100100001010010", 20293 => "1101000000001011", 20294 => "1001000011100001", 20295 => "1001001001000111", 20296 => "1101010111000100", 20297 => "1010111111100011", 20298 => "1110011010111101", 20299 => "0111101101011100", 20300 => "0001010011110010", 20301 => "0011111011000001", 20302 => "1010011101100101", 20303 => "0111011111000011", 20304 => "0111101001100011", 20305 => "1101101100101011", 20306 => "1000101011110111", 20307 => "1001011110011101", 20308 => "0001111010000001", 20309 => "1011000010111010", 20310 => "0000111001101011", 20311 => "0011001100111101", 20312 => "1111010110011111", 20313 => "1001111001000010", 20314 => "0111111001110100", 20315 => "0000101100100000", 20316 => "0110110010101001", 20317 => "1001100000100011", 20318 => "1101101011000011", 20319 => "1010111011001000", 20320 => "0001000101110011", 20321 => "1001110000000000", 20322 => "1010010101000010", 20323 => "0111100001110000", 20324 => "0100110100011100", 20325 => "0100000100111110", 20326 => "0100100111101000", 20327 => "0111110101100000", 20328 => "0000110101011100", 20329 => "0011110101110101", 20330 => "1111000110101101", 20331 => "0000110000010100", 20332 => "1010100110101000", 20333 => "0100010010101001", 20334 => "1001110111100001", 20335 => "1101010000101010", 20336 => "0110010011100011", 20337 => "0000011001110001", 20338 => "1010101100000111", 20339 => "1010100101110101", 20340 => "0100101100100101", 20341 => "1010001100111011", 20342 => "0111111100110100", 20343 => "0110110100110101", 20344 => "0010111000101100", 20345 => "0000010011000011", 20346 => "1111010011100111", 20347 => "0101100001011001", 20348 => "0110101011011011", 20349 => "1110000100001101", 20350 => "0110111100011101", 20351 => "0010111001001000", 20352 => "1101110101100011", 20353 => "1100101100101110", 20354 => "0100110001001010", 20355 => "1001001001100010", 20356 => "1101101111111110", 20357 => "0011100011011101", 20358 => "1001011111011001", 20359 => "0111111100001111", 20360 => "1000011000011001", 20361 => "1011011011111000", 20362 => "0110101111011110", 20363 => "1110110101010101", 20364 => "1101001100100011", 20365 => "1101111111001010", 20366 => "0101000011111000", 20367 => "0001101001100110", 20368 => "0001111111111001", 20369 => "0001110000010110", 20370 => "0101001101011011", 20371 => "1101110111011000", 20372 => "1101001001101000", 20373 => "0011111111011111", 20374 => "1011110010101101", 20375 => "1110111110101101", 20376 => "0111101010000011", 20377 => "0010111100110000", 20378 => "0101101001001111", 20379 => "1011101111100101", 20380 => "0001101010001000", 20381 => "0110011100100101", 20382 => "1001101101110101", 20383 => "0001110001001111", 20384 => "0000000010010100", 20385 => "1010010111001100", 20386 => "0010101111111010", 20387 => "0010100011010001", 20388 => "0011001010001001", 20389 => "1001100010010000", 20390 => "0010010000000111", 20391 => "1101000111011110", 20392 => "1111000011011011", 20393 => "0010110010010001", 20394 => "0011101000110010", 20395 => "1010001001001011", 20396 => "1111011000100011", 20397 => "1000001111010000", 20398 => "1010010101110010", 20399 => "1010010100110011", 20400 => "1001111110010011", 20401 => "1001101111000100", 20402 => "0011101100001101", 20403 => "1001110100100101", 20404 => "1111101101000001", 20405 => "0000100100101101", 20406 => "0010111011001011", 20407 => "1010111000010011", 20408 => "0000101011110101", 20409 => "0100000100111011", 20410 => "1100111011111110", 20411 => "1011000011001101", 20412 => "0110100000010000", 20413 => "0111000110101010", 20414 => "0011110100100100", 20415 => "0010010110101100", 20416 => "0110011011110111", 20417 => "1000011110010101", 20418 => "0001011011000011", 20419 => "1111010111011010", 20420 => "1100111011001100", 20421 => "0111101011100001", 20422 => "1111101000001001", 20423 => "0000000100100100", 20424 => "1001001101110111", 20425 => "0010101001010010", 20426 => "0011110010111011", 20427 => "1011111011110010", 20428 => "0101011111000101", 20429 => "1010111111010110", 20430 => "1010100011100010", 20431 => "1101111100001011", 20432 => "1000011000111100", 20433 => "1011110110011000", 20434 => "1000010001001001", 20435 => "1110100111000000", 20436 => "1010000101010000", 20437 => "0110001010110001", 20438 => "0000100110111001", 20439 => "1110011011101101", 20440 => "1110011101000111", 20441 => "0110110100101110", 20442 => "1000101111110111", 20443 => "0011011100000000", 20444 => "1100110110110000", 20445 => "0101000001011011", 20446 => "0100001010100101", 20447 => "1001100010110111", 20448 => "1101010000001111", 20449 => "0010000101000111", 20450 => "1100101011001011", 20451 => "1101111110111010", 20452 => "1000011010001111", 20453 => "0100111001101100", 20454 => "1111110110101110", 20455 => "0110101110100100", 20456 => "1000101011110010", 20457 => "0010010100010001", 20458 => "1010010001100010", 20459 => "0010101111001011", 20460 => "1010111000100111", 20461 => "0111010000101000", 20462 => "0000100001100111", 20463 => "0001110101101011", 20464 => "1100101100000101", 20465 => "0011110011011010", 20466 => "1101111011000000", 20467 => "1100010101001001", 20468 => "0101110011001111", 20469 => "0110111110000010", 20470 => "1011001000010011", 20471 => "0100001111101110", 20472 => "1110000100010110", 20473 => "0011011100111011", 20474 => "1101001010001101", 20475 => "0111100000101100", 20476 => "1110100000110100", 20477 => "1011000111000110", 20478 => "1100101101001010", 20479 => "0011000001110101", 20480 => "0010000111110111", 20481 => "0000101100110100", 20482 => "0101111101100010", 20483 => "1001010100001011", 20484 => "1000100010010110", 20485 => "0001101101101110", 20486 => "0100110101001000", 20487 => "0111111001111001", 20488 => "1111010010101000", 20489 => "1100000110000000", 20490 => "1010000100110100", 20491 => "0001010110011111", 20492 => "1000101010100111", 20493 => "0001111011111110", 20494 => "1001011110100100", 20495 => "1011001111111001", 20496 => "1101010101111111", 20497 => "1000011100100101", 20498 => "0010110110101010", 20499 => "0010110000101110", 20500 => "0001000001011011", 20501 => "0011110000101100", 20502 => "1010001011100010", 20503 => "0100110111001100", 20504 => "0010110101001111", 20505 => "1000110010110110", 20506 => "1111111101010001", 20507 => "1000001110010110", 20508 => "1111010011001010", 20509 => "0001101100010110", 20510 => "1100001110101101", 20511 => "1010100011011101", 20512 => "0110100010100010", 20513 => "1000010000100011", 20514 => "0010101110111001", 20515 => "0101101111111011", 20516 => "0001100101001010", 20517 => "0001111110011001", 20518 => "0100010011111011", 20519 => "1000000010100101", 20520 => "1000001011110110", 20521 => "0010101111111010", 20522 => "1000100111000000", 20523 => "0110110110010111", 20524 => "1110000101110101", 20525 => "0101010010011111", 20526 => "0010110111111001", 20527 => "1100100010001000", 20528 => "0110111111100111", 20529 => "1101110001101110", 20530 => "1101101100100100", 20531 => "1011010010101110", 20532 => "1111000111010101", 20533 => "0001110000001000", 20534 => "1110101101101111", 20535 => "1010000100010000", 20536 => "1110001110101011", 20537 => "0000011010001111", 20538 => "1100100010111010", 20539 => "1010111000010001", 20540 => "0011111100001000", 20541 => "1101011101011001", 20542 => "1001100011110110", 20543 => "0110010010110111", 20544 => "1000011100000100", 20545 => "1100000101111001", 20546 => "1000001110101100", 20547 => "1011111000100110", 20548 => "1110011111111000", 20549 => "0100101011101000", 20550 => "0111110101011011", 20551 => "0101100000100110", 20552 => "1110010111111000", 20553 => "1010110101000100", 20554 => "1101011011010110", 20555 => "1100111110101100", 20556 => "1110001110101110", 20557 => "0000000100011111", 20558 => "0111100100000110", 20559 => "0011011100011101", 20560 => "0001010010011111", 20561 => "1010111110011011", 20562 => "0011001111100000", 20563 => "0001110000011110", 20564 => "0100110101101000", 20565 => "1101111010011010", 20566 => "1001000101010111", 20567 => "1010011001101101", 20568 => "1000101011000011", 20569 => "0110110000001110", 20570 => "1001000010110010", 20571 => "0100110101000100", 20572 => "1000001101110011", 20573 => "1010110111100111", 20574 => "0000110010101000", 20575 => "1010100100110011", 20576 => "1111011101101000", 20577 => "0010000010100100", 20578 => "0110111010011001", 20579 => "0010000000111000", 20580 => "0011000000010110", 20581 => "1001001100001001", 20582 => "1110000111010111", 20583 => "0111101111100110", 20584 => "1001100001011011", 20585 => "1101110100101100", 20586 => "1100100110101011", 20587 => "0000001101100011", 20588 => "1011101110101100", 20589 => "1110000100001111", 20590 => "0111000001001000", 20591 => "1110110011110000", 20592 => "0111110101011101", 20593 => "1111011001011110", 20594 => "0000100100100100", 20595 => "1000101101111010", 20596 => "0101010010011110", 20597 => "1001010010011010", 20598 => "0111011011011001", 20599 => "0110011100110010", 20600 => "1011110000010101", 20601 => "0110001000101011", 20602 => "1100011000000111", 20603 => "0000010000011110", 20604 => "0000001110010110", 20605 => "0000010010011111", 20606 => "1100111100001100", 20607 => "0001110010011011", 20608 => "0100001100000101", 20609 => "0000000111110011", 20610 => "1100100110000011", 20611 => "1110111101110101", 20612 => "0100110011010000", 20613 => "0011001100010101", 20614 => "0011101000000110", 20615 => "0101010001011110", 20616 => "0101101110011011", 20617 => "0111010101101110", 20618 => "0100100010111101", 20619 => "1101011100000000", 20620 => "1110111100001000", 20621 => "0010101111011100", 20622 => "0000101011010111", 20623 => "1001101111100010", 20624 => "1110000110000010", 20625 => "1001001100010100", 20626 => "0110000100000010", 20627 => "1101101010110011", 20628 => "0101110000101111", 20629 => "1011001101011100", 20630 => "0010001000111010", 20631 => "1101111011010101", 20632 => "0011100101111110", 20633 => "1011001011010010", 20634 => "0111110110111000", 20635 => "1111101110110101", 20636 => "1011110111001011", 20637 => "0110101000111100", 20638 => "0010100101111100", 20639 => "1111000110110101", 20640 => "1101100011100100", 20641 => "1011011011000011", 20642 => "1110111100101110", 20643 => "1100101111100110", 20644 => "1011001110111000", 20645 => "0101101110110011", 20646 => "1011000000100000", 20647 => "1111110001010010", 20648 => "0010101001011000", 20649 => "0111100001001101", 20650 => "1100111101010011", 20651 => "0101011011011011", 20652 => "1111110000010001", 20653 => "0001110100001000", 20654 => "1111011011101100", 20655 => "1111001001111001", 20656 => "1101111001101100", 20657 => "0101011000000000", 20658 => "1011011101100111", 20659 => "1110100111010101", 20660 => "0111101101010000", 20661 => "1101110001101111", 20662 => "0111010100001110", 20663 => "0100010110010000", 20664 => "0101111111011001", 20665 => "0101000001011101", 20666 => "1111000011100001", 20667 => "1011000000010011", 20668 => "1010010110001010", 20669 => "0101010110001001", 20670 => "0001001001001010", 20671 => "0000111000011100", 20672 => "0001001100011010", 20673 => "1010110101111011", 20674 => "1101101110110000", 20675 => "1000101110100010", 20676 => "1101101111100010", 20677 => "0001000110000101", 20678 => "1001101001100100", 20679 => "0101011000001100", 20680 => "0010011111001001", 20681 => "1111100001000100", 20682 => "0110101110111101", 20683 => "1010101100101101", 20684 => "1001100101101101", 20685 => "1110001100000101", 20686 => "0001110100000010", 20687 => "0101101011110000", 20688 => "0000110101110111", 20689 => "1010011101110100", 20690 => "1110000100101000", 20691 => "1111000111110100", 20692 => "0010010000111101", 20693 => "1111010011000001", 20694 => "0000100000000101", 20695 => "1101010110110010", 20696 => "1110101111001000", 20697 => "0010000111101000", 20698 => "1010111000001000", 20699 => "1000101110101001", 20700 => "1110010011111111", 20701 => "0111001101110011", 20702 => "0111000001100011", 20703 => "1000001011000010", 20704 => "0110101111101110", 20705 => "1101100001000100", 20706 => "1011000010100010", 20707 => "1101100010101001", 20708 => "0001100110000001", 20709 => "1110011111101010", 20710 => "0000110100010110", 20711 => "0100110001111110", 20712 => "0111110010100001", 20713 => "1111101101101001", 20714 => "1011111110001101", 20715 => "1100111001111101", 20716 => "1001001000100000", 20717 => "1111010000101010", 20718 => "0100000110000010", 20719 => "0001010010111001", 20720 => "0011101000010000", 20721 => "0000011111001110", 20722 => "0001111111010011", 20723 => "1110010110001011", 20724 => "1010011101100111", 20725 => "1001011100110010", 20726 => "0111010111110010", 20727 => "0100100110111011", 20728 => "1100010101011001", 20729 => "1011110110100100", 20730 => "0001011101011011", 20731 => "0000000101000100", 20732 => "1100110001101000", 20733 => "0101111110100000", 20734 => "0100111011010001", 20735 => "0001111100010010", 20736 => "1001010100001001", 20737 => "0101000011010001", 20738 => "0100100101000000", 20739 => "0011001111010001", 20740 => "0110001011010100", 20741 => "0110001100011110", 20742 => "0111011100011010", 20743 => "1110111011000111", 20744 => "0000100011011000", 20745 => "1000000001011010", 20746 => "0011110111110000", 20747 => "1111111001000101", 20748 => "0111000010010110", 20749 => "0110110011100111", 20750 => "1001111001110100", 20751 => "1011011000100011", 20752 => "1110111000010011", 20753 => "0001000100000011", 20754 => "0001101000111100", 20755 => "1101000101110110", 20756 => "0000110100000001", 20757 => "1110100010000101", 20758 => "0100110011101110", 20759 => "0010110011101111", 20760 => "0000011111001001", 20761 => "0010000001001000", 20762 => "0101110001110001", 20763 => "1000101000000101", 20764 => "0101010010100110", 20765 => "0010101111111110", 20766 => "0100001001000001", 20767 => "1110001100110101", 20768 => "0000011110110101", 20769 => "0111011100100000", 20770 => "0111100000110100", 20771 => "0110101110011110", 20772 => "1100100100100110", 20773 => "0000110000001101", 20774 => "0011010000000000", 20775 => "1111111111011111", 20776 => "1111101001100011", 20777 => "1011010011110111", 20778 => "0010001010001110", 20779 => "0100011000100100", 20780 => "1101010010110010", 20781 => "0101010001100011", 20782 => "1000010001110110", 20783 => "0100011111000100", 20784 => "0101101011011001", 20785 => "0001111011011000", 20786 => "0000111111001010", 20787 => "1001100010011111", 20788 => "0110111100110100", 20789 => "1011101101001010", 20790 => "0100001100010000", 20791 => "0111000111111000", 20792 => "0001111000000011", 20793 => "1010010001111111", 20794 => "1011110101001111", 20795 => "1000001000001000", 20796 => "1101001000101011", 20797 => "0000101111100010", 20798 => "1110010000001000", 20799 => "0110100111011100", 20800 => "1111111100010111", 20801 => "1011001010001001", 20802 => "1111100101010001", 20803 => "1111100111010010", 20804 => "1011001110010001", 20805 => "0010110110101111", 20806 => "1000110000011100", 20807 => "0001001000001000", 20808 => "1001010100110110", 20809 => "1110011001100111", 20810 => "1110110000111011", 20811 => "1001100011100101", 20812 => "0010100111011011", 20813 => "1111100100111100", 20814 => "0010110101100100", 20815 => "0011100100011100", 20816 => "0000000001010101", 20817 => "1110000111101010", 20818 => "0100001111011001", 20819 => "1011001001010001", 20820 => "0010111110010110", 20821 => "1011110100111100", 20822 => "0111001010110011", 20823 => "1010000010001011", 20824 => "0101011000100011", 20825 => "0001110010100010", 20826 => "0000010001100111", 20827 => "1010101000111000", 20828 => "1010111111111000", 20829 => "1100111100001111", 20830 => "0000010010101101", 20831 => "0101011100011110", 20832 => "0010011101110001", 20833 => "1010001010111111", 20834 => "1111000000000110", 20835 => "1110100001100011", 20836 => "1001110011100101", 20837 => "1110000101111011", 20838 => "1001001100111001", 20839 => "0100001000101101", 20840 => "1100111111000001", 20841 => "0111101000100011", 20842 => "1101000010110111", 20843 => "0001100001101100", 20844 => "1000011111110001", 20845 => "1011110010101001", 20846 => "1010110101111111", 20847 => "1000111101100000", 20848 => "0000010001101100", 20849 => "1110001111010101", 20850 => "0010111010010000", 20851 => "0110001100111011", 20852 => "0101000110011101", 20853 => "0001110000000001", 20854 => "0000111101011111", 20855 => "0000001001000101", 20856 => "0011000101000100", 20857 => "0111010111011001", 20858 => "0100001110100101", 20859 => "0110111001111110", 20860 => "1111100111100110", 20861 => "0110001111101110", 20862 => "0100001100010011", 20863 => "0110110001000000", 20864 => "1000011100010100", 20865 => "1111011011010100", 20866 => "0100101000010010", 20867 => "1000110010110101", 20868 => "1000011110110110", 20869 => "0111110110101000", 20870 => "0011000111001101", 20871 => "1011001111001110", 20872 => "1111101011010110", 20873 => "0111000110011010", 20874 => "1100000110100110", 20875 => "0100110000110011", 20876 => "1111000110001011", 20877 => "0111110001000011", 20878 => "1100110100101000", 20879 => "1111100101100011", 20880 => "1000011011000110", 20881 => "1101011100110100", 20882 => "1100011010100100", 20883 => "1110101010000101", 20884 => "1001000001110010", 20885 => "1101111111100001", 20886 => "1001110011101111", 20887 => "1111110000110010", 20888 => "1110000101110010", 20889 => "0000000000111010", 20890 => "1100011110100001", 20891 => "1010111110110111", 20892 => "1010010000100000", 20893 => "1101111001001000", 20894 => "0001110110010111", 20895 => "0000011011011001", 20896 => "1111010110010101", 20897 => "0111010110001011", 20898 => "0101110110001101", 20899 => "1000101100100000", 20900 => "1100011100101010", 20901 => "1111000101100101", 20902 => "0001010101010010", 20903 => "0010000100101101", 20904 => "0110101111001101", 20905 => "0101110110000110", 20906 => "1010001011111110", 20907 => "1001000111000010", 20908 => "1110100010001100", 20909 => "0100010011110001", 20910 => "0110010100110000", 20911 => "0110110110010110", 20912 => "1011111000101001", 20913 => "0100110101101010", 20914 => "1101101101000000", 20915 => "1010001000110010", 20916 => "1010111010000111", 20917 => "1011110111001100", 20918 => "1000110001011000", 20919 => "0000100011111010", 20920 => "1011111100110011", 20921 => "0111100111111111", 20922 => "0111011011101010", 20923 => "1101110011100001", 20924 => "1101110101100001", 20925 => "1010100001101100", 20926 => "1010010101000001", 20927 => "0111101110011101", 20928 => "1110101110111001", 20929 => "0010011000000101", 20930 => "1001010111010000", 20931 => "1000001000000000", 20932 => "0011010110001100", 20933 => "0111101101000110", 20934 => "1110111111010000", 20935 => "0110011011110100", 20936 => "0100101011010010", 20937 => "1100011010101111", 20938 => "0111110100000011", 20939 => "0010111111001110", 20940 => "1010110111111110", 20941 => "0101001110100010", 20942 => "0100001001101001", 20943 => "0110001111000011", 20944 => "1101111110100110", 20945 => "1000100100111010", 20946 => "1011111000011101", 20947 => "0000110000110101", 20948 => "0011010001000010", 20949 => "0101000101111000", 20950 => "0000000010101001", 20951 => "0011010110000011", 20952 => "0100000100011011", 20953 => "1011000101100000", 20954 => "1110110011100000", 20955 => "1111101100010000", 20956 => "0101010011110000", 20957 => "0001101110100001", 20958 => "0110011011011011", 20959 => "1101110001100010", 20960 => "1011100001100001", 20961 => "0101111011001001", 20962 => "1101101011111001", 20963 => "1000111011001101", 20964 => "1110110111001111", 20965 => "0101111010110110", 20966 => "1000100110011011", 20967 => "0111100010011111", 20968 => "0100111010001111", 20969 => "0011011010011110", 20970 => "1001111110010010", 20971 => "0000010110110111", 20972 => "0110110010001010", 20973 => "1010100001100001", 20974 => "1100110000011011", 20975 => "1101011100110110", 20976 => "1011111001111001", 20977 => "1011010010010000", 20978 => "1110011110010001", 20979 => "1101101100011111", 20980 => "1100010111011100", 20981 => "0100010011111000", 20982 => "0011110000010011", 20983 => "0011011111111001", 20984 => "1001110100111000", 20985 => "1011100110000100", 20986 => "0001011001110001", 20987 => "0001010001000010", 20988 => "0010000101000010", 20989 => "0110000010011100", 20990 => "0101011111101010", 20991 => "1000101100101100", 20992 => "0101110001101111", 20993 => "1101101011010010", 20994 => "0001101110010101", 20995 => "0100011100110001", 20996 => "0101001101011100", 20997 => "1000100010111000", 20998 => "1001110000101111", 20999 => "0101000111100110", 21000 => "1000001100100101", 21001 => "0000110100100010", 21002 => "0010011111100101", 21003 => "0010011011010111", 21004 => "0011100010010010", 21005 => "0100010101110111", 21006 => "0101111111111001", 21007 => "1111110001010100", 21008 => "0011001111100110", 21009 => "1100101000001010", 21010 => "0011110000000000", 21011 => "1110001010100000", 21012 => "1101001111001011", 21013 => "0001101111000000", 21014 => "0100000011001001", 21015 => "1111111110000111", 21016 => "0101111001010010", 21017 => "1101000010001111", 21018 => "1100101101011110", 21019 => "0101100110011101", 21020 => "1111111101101110", 21021 => "0100001110010111", 21022 => "1100100010010010", 21023 => "1000000011101001", 21024 => "0101101010111000", 21025 => "0011010111001101", 21026 => "0010010111100111", 21027 => "0101000111010101", 21028 => "1111011001101110", 21029 => "1000100000101001", 21030 => "1101010000101110", 21031 => "1000001111111000", 21032 => "0010011110010001", 21033 => "1000100000010001", 21034 => "0100010110110101", 21035 => "0000100111110011", 21036 => "0100111011101001", 21037 => "1101111011011101", 21038 => "1101000111110000", 21039 => "0000100100001100", 21040 => "0000110111010001", 21041 => "1110111011110010", 21042 => "0010011101101000", 21043 => "0010000011111011", 21044 => "0100011101110001", 21045 => "1111011000100001", 21046 => "1111110111110101", 21047 => "1101111000010111", 21048 => "0000111101010001", 21049 => "0100011111111110", 21050 => "1011001010110101", 21051 => "1010001000010000", 21052 => "1110000000100100", 21053 => "1011110101111010", 21054 => "1011100011000110", 21055 => "0101001110100001", 21056 => "1001001110101010", 21057 => "1101001001010101", 21058 => "0010010010011100", 21059 => "0100010110001100", 21060 => "0010000100011110", 21061 => "1111010001000010", 21062 => "1101010010111101", 21063 => "0001001011010111", 21064 => "0111011101011100", 21065 => "0011111111011101", 21066 => "1110111110101010", 21067 => "1100000101011101", 21068 => "1111010110000011", 21069 => "1100110001100001", 21070 => "1110000111010000", 21071 => "0011010011110101", 21072 => "1011010011100101", 21073 => "0000110110000100", 21074 => "1011000010001011", 21075 => "1100000110111001", 21076 => "1011111010001111", 21077 => "0010011110000000", 21078 => "0100011100111110", 21079 => "0111000111100111", 21080 => "0001111000011011", 21081 => "0001010011101100", 21082 => "1011100110001101", 21083 => "1000101001101011", 21084 => "0101100101101000", 21085 => "1000011000101010", 21086 => "1111000110001111", 21087 => "0000010000001100", 21088 => "1000111100101010", 21089 => "0111011010100111", 21090 => "0011000011000111", 21091 => "0000010001010001", 21092 => "0101111110111100", 21093 => "1111010000110100", 21094 => "1111100111111000", 21095 => "0011110100101100", 21096 => "1010101000111000", 21097 => "1001100110001000", 21098 => "0001000011001001", 21099 => "1101001110010001", 21100 => "1001011011001011", 21101 => "0101000011101000", 21102 => "1101111110110100", 21103 => "0010110111011001", 21104 => "1110001111100111", 21105 => "0011011011010001", 21106 => "1111110000000100", 21107 => "0110000010011000", 21108 => "0110001111010111", 21109 => "1101000111010110", 21110 => "0000011101010110", 21111 => "0100110101000011", 21112 => "0001111000110101", 21113 => "1101001001101010", 21114 => "1010000110010010", 21115 => "1101010111101000", 21116 => "0111110110010100", 21117 => "0000011000101110", 21118 => "1100101010010000", 21119 => "0000100111010000", 21120 => "0010001001001111", 21121 => "1010101010100111", 21122 => "0101010111110010", 21123 => "0001001010000110", 21124 => "1011001010110111", 21125 => "1100010111000011", 21126 => "0001110000100010", 21127 => "1001111010100010", 21128 => "0000001001010111", 21129 => "0001110001100101", 21130 => "0010111010111101", 21131 => "0000111010010001", 21132 => "1101111111010110", 21133 => "0001000010010100", 21134 => "1011110000101100", 21135 => "0001010101001001", 21136 => "0111101000110010", 21137 => "1000111110000011", 21138 => "1100111011110010", 21139 => "0011001000011101", 21140 => "1011111110100000", 21141 => "0010001010011001", 21142 => "1001000100111110", 21143 => "0010011010100100", 21144 => "0111111001011111", 21145 => "0110110010010100", 21146 => "1011101000110100", 21147 => "1001101010000011", 21148 => "0000110111011000", 21149 => "0011011111000010", 21150 => "1100001010001111", 21151 => "0110100100110100", 21152 => "1001010101010101", 21153 => "0000111100010000", 21154 => "0110011101010100", 21155 => "0111111000111111", 21156 => "1101101110100100", 21157 => "0110010101010011", 21158 => "0100110001011101", 21159 => "1010100000001011", 21160 => "0001110001000110", 21161 => "1010011011001110", 21162 => "0010111010011100", 21163 => "0011001011101001", 21164 => "0000001100101111", 21165 => "0010110111101110", 21166 => "1001111010101010", 21167 => "1100001010110111", 21168 => "0000011111011010", 21169 => "1000011100100100", 21170 => "1111110100101000", 21171 => "1110001110101001", 21172 => "0001010101111100", 21173 => "1110010111101100", 21174 => "0011000101100110", 21175 => "1111101010001000", 21176 => "1100110100110100", 21177 => "0011111101111101", 21178 => "1001110001101110", 21179 => "1011010110110010", 21180 => "1000010010010101", 21181 => "1110000101010011", 21182 => "1011101010100100", 21183 => "1100000101111110", 21184 => "0111001110101001", 21185 => "0110111011011101", 21186 => "0111000101010111", 21187 => "1111010100001100", 21188 => "1100000100100110", 21189 => "1000101101110101", 21190 => "1111010111000001", 21191 => "1100001010101000", 21192 => "1000010001100001", 21193 => "1010011001011100", 21194 => "1000111000100011", 21195 => "0000100001111011", 21196 => "1100001101101111", 21197 => "0100101110100001", 21198 => "1001101000100010", 21199 => "1110011010111110", 21200 => "1011101110010011", 21201 => "1100011000101101", 21202 => "1100001110110001", 21203 => "1101110001001011", 21204 => "1000010001110110", 21205 => "1001101011100000", 21206 => "1010110001001110", 21207 => "0100010110110010", 21208 => "0101110010111000", 21209 => "0101010100011111", 21210 => "0110101110110100", 21211 => "0101000100101100", 21212 => "0100110001011110", 21213 => "0110011111011011", 21214 => "1100110011101111", 21215 => "1001111101001101", 21216 => "0101011100011101", 21217 => "1000011111001110", 21218 => "1001000011101111", 21219 => "1110101100101101", 21220 => "0111010010110100", 21221 => "1100001100001110", 21222 => "1010110111010100", 21223 => "1000101011111111", 21224 => "0010001111111011", 21225 => "1101110000101101", 21226 => "0010101100000000", 21227 => "0110111000001110", 21228 => "0011100100001001", 21229 => "0011110000010011", 21230 => "1100111100010111", 21231 => "1000010111000010", 21232 => "0110011010000011", 21233 => "1110011001101110", 21234 => "1101100010111111", 21235 => "1111001111011101", 21236 => "1111010001011010", 21237 => "1111110001011000", 21238 => "0010000111111101", 21239 => "0010101111111001", 21240 => "0000011011011110", 21241 => "0100110100110001", 21242 => "0000001011100011", 21243 => "0000111010110101", 21244 => "1111101111110110", 21245 => "1010111101011010", 21246 => "0110101110111001", 21247 => "0001011001111111", 21248 => "0110100010101100", 21249 => "0111100011110101", 21250 => "1000011010110001", 21251 => "0111000011001011", 21252 => "1111010111010100", 21253 => "1100010100100011", 21254 => "0001011000001010", 21255 => "1101010010110100", 21256 => "0000010010001001", 21257 => "1011110000001000", 21258 => "0111111010010101", 21259 => "0010010000100000", 21260 => "1001000001000110", 21261 => "0010010111011001", 21262 => "1000011001001001", 21263 => "0000011000010001", 21264 => "0100000010101010", 21265 => "1011111110011001", 21266 => "0011011111110111", 21267 => "0010010101011110", 21268 => "0110111001010110", 21269 => "1000001001111010", 21270 => "0101011000000001", 21271 => "0110000011100111", 21272 => "1110010110110101", 21273 => "1111111010011110", 21274 => "1100011010100111", 21275 => "0001010011111000", 21276 => "1011000010001111", 21277 => "1010100010100110", 21278 => "1100111001110101", 21279 => "0000001010101100", 21280 => "0011110001110110", 21281 => "0001011101001001", 21282 => "1010101011010111", 21283 => "0101000011010011", 21284 => "0110110110001101", 21285 => "1011101101010100", 21286 => "0100001111101100", 21287 => "1110110100001011", 21288 => "0011011000011001", 21289 => "0011010000000111", 21290 => "1011110111001100", 21291 => "1001100101000110", 21292 => "0100101100010110", 21293 => "1111001001000110", 21294 => "1000101000001101", 21295 => "1100110101001110", 21296 => "0110001110111010", 21297 => "0001100110110011", 21298 => "0111011001011111", 21299 => "0110011101100001", 21300 => "1110100111000000", 21301 => "1100000100001111", 21302 => "1101111000011110", 21303 => "0110110111000001", 21304 => "1111000100001111", 21305 => "0011110010010100", 21306 => "0010111100001010", 21307 => "0000000001001010", 21308 => "1010001110110001", 21309 => "0001001110000110", 21310 => "0101011100100011", 21311 => "0011101011011100", 21312 => "1001101110101111", 21313 => "1100110010110101", 21314 => "1011101001101111", 21315 => "1010110001100000", 21316 => "1010110011111001", 21317 => "0110101110101101", 21318 => "1000101111000111", 21319 => "0110000001000111", 21320 => "1011111001111000", 21321 => "1001000101111101", 21322 => "0111101100100000", 21323 => "1111010110000100", 21324 => "0010110100101000", 21325 => "0010000110110100", 21326 => "0010111111101101", 21327 => "1101001110000011", 21328 => "1000111100110101", 21329 => "1010011101111011", 21330 => "1100011000110001", 21331 => "1000111101110100", 21332 => "1010001111110001", 21333 => "1000111000111101", 21334 => "1101010101000000", 21335 => "1110000101010111", 21336 => "1011011011110000", 21337 => "0100110000000101", 21338 => "0011000000001101", 21339 => "0111001101100011", 21340 => "0000111001000100", 21341 => "1111011101110010", 21342 => "0001011011001101", 21343 => "1000010111100001", 21344 => "1011100100001000", 21345 => "0100110111100111", 21346 => "1000010110101110", 21347 => "1000010100111000", 21348 => "0111110111011110", 21349 => "0011000101101010", 21350 => "1110110100001011", 21351 => "1011111010100000", 21352 => "1001010010000101", 21353 => "1110100000101111", 21354 => "1100101101111110", 21355 => "0010000110000110", 21356 => "1101011000010010", 21357 => "1110000000010010", 21358 => "0100100111101000", 21359 => "1001001101011000", 21360 => "0101011111101110", 21361 => "0011110101001100", 21362 => "1000111101001010", 21363 => "1111000111110000", 21364 => "1111101100110000", 21365 => "1010111101110000", 21366 => "0100000110110101", 21367 => "0110111100101101", 21368 => "1000001000111000", 21369 => "0110000010011011", 21370 => "0100110010101101", 21371 => "1110010001010000", 21372 => "1011001001101101", 21373 => "1011110100110100", 21374 => "0000100000100010", 21375 => "1110110000101011", 21376 => "0001001011011011", 21377 => "1011001110110111", 21378 => "0010011110110111", 21379 => "0000100110011011", 21380 => "1101000100000111", 21381 => "1000011110001011", 21382 => "1101110001010000", 21383 => "0011101000000100", 21384 => "1100001100010111", 21385 => "0111001110000111", 21386 => "0101010100010001", 21387 => "0010000001001100", 21388 => "1010100000100101", 21389 => "1110111010001001", 21390 => "1000100011000001", 21391 => "1110000100001001", 21392 => "0100000001010110", 21393 => "1110111100011111", 21394 => "0101001111000011", 21395 => "1111001101001101", 21396 => "0000110010010101", 21397 => "1101100011101000", 21398 => "1110010100001010", 21399 => "0100010011011001", 21400 => "1101101010111001", 21401 => "0111110011100011", 21402 => "1010101101101001", 21403 => "0011111110000010", 21404 => "0111010110111100", 21405 => "1110110110111100", 21406 => "0111110100001111", 21407 => "1111100111000001", 21408 => "0101100110111110", 21409 => "1110000100111100", 21410 => "1100100100000101", 21411 => "1010000100100101", 21412 => "0011110111100110", 21413 => "0101000011001110", 21414 => "1110011111010100", 21415 => "0011110000110001", 21416 => "1010011001001001", 21417 => "0110111011100111", 21418 => "1100100011011101", 21419 => "0010110001100110", 21420 => "0001001110011100", 21421 => "0010010100000110", 21422 => "1100101010001111", 21423 => "1000100000101111", 21424 => "0101110100000010", 21425 => "0111011100001011", 21426 => "1110100111000111", 21427 => "0010101011010011", 21428 => "0111010100000010", 21429 => "0100101011000101", 21430 => "0110100010011000", 21431 => "1100001110010010", 21432 => "1010101011101000", 21433 => "0000010000100100", 21434 => "0111101100100111", 21435 => "1001011101110100", 21436 => "1000101011000110", 21437 => "0011001110011100", 21438 => "0011010110101000", 21439 => "1011111110010111", 21440 => "1101100011001101", 21441 => "0110001010100010", 21442 => "0010100101111001", 21443 => "1011111111110100", 21444 => "1011110110111110", 21445 => "0010111011100100", 21446 => "0011101011001110", 21447 => "1000010001000101", 21448 => "0000100110001111", 21449 => "0101110000100101", 21450 => "0011111000010000", 21451 => "0000000110101101", 21452 => "0011110111101011", 21453 => "1101101011010001", 21454 => "0000010111110001", 21455 => "0001010100101110", 21456 => "1101101111101111", 21457 => "0000010010001100", 21458 => "0110010001111001", 21459 => "0110111010110110", 21460 => "1100110101010110", 21461 => "0111111001011110", 21462 => "0010101111111101", 21463 => "1011100011010101", 21464 => "0100101110100001", 21465 => "1000001010001111", 21466 => "1110010011000100", 21467 => "1110111000011011", 21468 => "1001100100100110", 21469 => "0101010001110001", 21470 => "0001001111110011", 21471 => "0110101100100100", 21472 => "0001000010101010", 21473 => "0100110001011101", 21474 => "0110000111111001", 21475 => "0110011100010100", 21476 => "1011100000001110", 21477 => "1011111010101110", 21478 => "0100100100001110", 21479 => "1110111001111101", 21480 => "0111001001110011", 21481 => "0101010000100101", 21482 => "0111001101000010", 21483 => "1110001110001001", 21484 => "0001111100110111", 21485 => "1000100110010000", 21486 => "1011110111110100", 21487 => "0101101101101011", 21488 => "1010010001111100", 21489 => "0000110110011011", 21490 => "1011101111000110", 21491 => "1011111010101111", 21492 => "0000111101101101", 21493 => "1000110100001110", 21494 => "1100011010010101", 21495 => "0001111010111110", 21496 => "1101010000010101", 21497 => "1000001111101111", 21498 => "0001100011100011", 21499 => "1000011000001100", 21500 => "0010111001101111", 21501 => "0111101110000100", 21502 => "0101011110100100", 21503 => "1010001111111001", 21504 => "1010100100001100", 21505 => "0011000010110000", 21506 => "1010010110101000", 21507 => "0100100101101111", 21508 => "0011011000101000", 21509 => "1010010110001000", 21510 => "0100111101001100", 21511 => "0100110000011111", 21512 => "0101110010100110", 21513 => "0100010000111011", 21514 => "1111001100110010", 21515 => "0010100001110010", 21516 => "1111011011011001", 21517 => "0011001101000110", 21518 => "1111000110110010", 21519 => "0000001110101010", 21520 => "1101110010110010", 21521 => "0010111101101010", 21522 => "1001101110100110", 21523 => "0101011001000010", 21524 => "1101110110111010", 21525 => "1100010011101011", 21526 => "1100001111010011", 21527 => "0001100110001100", 21528 => "1010010111100110", 21529 => "1011010100001100", 21530 => "0000100011111010", 21531 => "1100101000001001", 21532 => "1111101101110101", 21533 => "0011100000100000", 21534 => "0110000010010010", 21535 => "0010001001110110", 21536 => "1001111100001100", 21537 => "0000011111111011", 21538 => "1100100100000101", 21539 => "1000010110111110", 21540 => "1001101110010001", 21541 => "1000010011010010", 21542 => "1101111001111000", 21543 => "0011010101001010", 21544 => "1101010000110111", 21545 => "1101011110111010", 21546 => "1100101011111111", 21547 => "1010011010011001", 21548 => "0001111111100100", 21549 => "0110000000101011", 21550 => "0100010111111000", 21551 => "1010110100010100", 21552 => "1011011101011101", 21553 => "1011001101111011", 21554 => "0101110110110111", 21555 => "1011110110100111", 21556 => "0001100001110001", 21557 => "0110011110010011", 21558 => "0100000111100010", 21559 => "1000011001010111", 21560 => "0110111100011100", 21561 => "1100001111110010", 21562 => "0010101100011100", 21563 => "1110110001111100", 21564 => "0110111011100101", 21565 => "1111011111111111", 21566 => "0101000011010011", 21567 => "1001011101010111", 21568 => "1110000000101011", 21569 => "0000011100101011", 21570 => "1000010001011110", 21571 => "1001011110110000", 21572 => "1100101000000100", 21573 => "1000100011001100", 21574 => "1000111010011101", 21575 => "0100001111011111", 21576 => "1010000011101101", 21577 => "0100010011011011", 21578 => "1011011100110000", 21579 => "1111110001010100", 21580 => "1000000001111101", 21581 => "0100011001011001", 21582 => "0001110000010111", 21583 => "1111101111011101", 21584 => "1100100000001111", 21585 => "0110110001110010", 21586 => "1111111001000011", 21587 => "1100101101101010", 21588 => "1101001011001100", 21589 => "0001000100011110", 21590 => "0001110010000100", 21591 => "0110101110111111", 21592 => "0110110010111001", 21593 => "0001001101111101", 21594 => "1110100010011100", 21595 => "1101110110100011", 21596 => "0000001111110111", 21597 => "1000001110000001", 21598 => "0100010110111111", 21599 => "0010100111101111", 21600 => "0100101100000010", 21601 => "0001000101001011", 21602 => "1000000000111001", 21603 => "0101100110010010", 21604 => "0000001100101001", 21605 => "0101111011000011", 21606 => "0111011111100100", 21607 => "0100001001111110", 21608 => "0100100011100110", 21609 => "0101101110001000", 21610 => "0100111000100110", 21611 => "0110000001100011", 21612 => "1001110011010010", 21613 => "1000101110010100", 21614 => "1100110101110000", 21615 => "0000010110011100", 21616 => "0110111100110110", 21617 => "0110101110100000", 21618 => "0001000110110010", 21619 => "1101101010000000", 21620 => "1000110101100011", 21621 => "0011011001110011", 21622 => "0110110110110101", 21623 => "1011000101101000", 21624 => "0001001010000010", 21625 => "0110101000110100", 21626 => "0101000101010110", 21627 => "1000111001101101", 21628 => "0011101110011001", 21629 => "1110000010100010", 21630 => "1001100000111010", 21631 => "0100111100001001", 21632 => "1000111000010110", 21633 => "1010000010011010", 21634 => "1000000001010010", 21635 => "1111011110011100", 21636 => "0110010000001100", 21637 => "0010010011011000", 21638 => "0010000000101110", 21639 => "0011011100010000", 21640 => "0100000111100000", 21641 => "1010100010001001", 21642 => "1111110001011100", 21643 => "0011110110100001", 21644 => "0101101010101100", 21645 => "0111000100100000", 21646 => "1001011010101101", 21647 => "1100110001001101", 21648 => "1000011000010000", 21649 => "0101100101001011", 21650 => "0001001011111110", 21651 => "0000000000101111", 21652 => "0101111111001011", 21653 => "0100001000000011", 21654 => "1111110101101110", 21655 => "1011000111011101", 21656 => "0000010111101011", 21657 => "0100100000101111", 21658 => "1111110011110100", 21659 => "0111010110000110", 21660 => "0011111001010111", 21661 => "1001011001111100", 21662 => "1101111011100011", 21663 => "1000011001010011", 21664 => "0110100000111100", 21665 => "1000110011001010", 21666 => "0010100100011101", 21667 => "1010101111100011", 21668 => "0111100110011110", 21669 => "1001010011100101", 21670 => "0010110110101100", 21671 => "0000011000011001", 21672 => "1101111010001101", 21673 => "0100110100001111", 21674 => "0111010111101001", 21675 => "1010001110001010", 21676 => "1110010010110111", 21677 => "1011010111111100", 21678 => "0101010000101010", 21679 => "1101101101010110", 21680 => "1100010110000111", 21681 => "1101001101000000", 21682 => "0101000110011110", 21683 => "1010100011000110", 21684 => "0001101000011001", 21685 => "1010111010010000", 21686 => "0110011111110000", 21687 => "1101100100010001", 21688 => "1001111111111111", 21689 => "0100001110111011", 21690 => "1000001110001110", 21691 => "1000011100000100", 21692 => "0011011000000010", 21693 => "0001111110100000", 21694 => "1101111000100101", 21695 => "0100110100101010", 21696 => "0111111100100100", 21697 => "0101001010111101", 21698 => "0101111010110100", 21699 => "1100000000000011", 21700 => "0110010001011110", 21701 => "1010110000101101", 21702 => "1000001111110001", 21703 => "1110001111011001", 21704 => "0010000110000110", 21705 => "0111100000110001", 21706 => "0000100100001111", 21707 => "1010111110011100", 21708 => "1101000010100100", 21709 => "0101100010001111", 21710 => "0010000011010000", 21711 => "0100100101110101", 21712 => "0000100010001011", 21713 => "0011111001101100", 21714 => "0101011100010111", 21715 => "0100010101110110", 21716 => "1010011111001101", 21717 => "1001011100111010", 21718 => "0001011001000100", 21719 => "0110001100110000", 21720 => "0001010110111000", 21721 => "0000111000011010", 21722 => "1101101101110111", 21723 => "0110101100001001", 21724 => "1001111111111100", 21725 => "1100000111011001", 21726 => "1101101111000110", 21727 => "0111100111001111", 21728 => "1111101001001010", 21729 => "1110101000011010", 21730 => "1010000011011010", 21731 => "1100100000101101", 21732 => "0100000111010011", 21733 => "1101011110001111", 21734 => "1111000111101001", 21735 => "0000000111011111", 21736 => "1111001000000000", 21737 => "1101001100011010", 21738 => "0110100000100110", 21739 => "1001110101001011", 21740 => "0001001110110010", 21741 => "1110101000001010", 21742 => "0110010000100111", 21743 => "0110110011010101", 21744 => "1001010100010101", 21745 => "1100000000000001", 21746 => "0011010101010100", 21747 => "0110111111101101", 21748 => "1111111011011110", 21749 => "1110110111110110", 21750 => "0000111001010101", 21751 => "1001110001100110", 21752 => "0001010001001000", 21753 => "1100100110000001", 21754 => "1111111011010110", 21755 => "1000111100001001", 21756 => "1011110100110010", 21757 => "0110101010110111", 21758 => "1010011011001111", 21759 => "0111010101100001", 21760 => "1010111001111111", 21761 => "0110110110000101", 21762 => "1000110100100110", 21763 => "1110111101100010", 21764 => "0111010001101010", 21765 => "0010100110010011", 21766 => "0111110111101100", 21767 => "0101110011110101", 21768 => "0000011101110000", 21769 => "1000101011111110", 21770 => "1110110100011101", 21771 => "0111101010000101", 21772 => "0011100010011001", 21773 => "0110110000110110", 21774 => "1000110000110101", 21775 => "0000000111110101", 21776 => "0011000100010001", 21777 => "0011011001001110", 21778 => "0110111010000011", 21779 => "1011100011100100", 21780 => "1010001110000101", 21781 => "0000110010111110", 21782 => "1100000000011001", 21783 => "1011011010011101", 21784 => "0100000010001110", 21785 => "1001110101001111", 21786 => "1101011110100011", 21787 => "1001000111010100", 21788 => "1001111111000111", 21789 => "0111011000010001", 21790 => "0111111001000111", 21791 => "1010000010110000", 21792 => "1000011101011110", 21793 => "1110110011010101", 21794 => "0010000111010110", 21795 => "0100101011010100", 21796 => "1000101001001100", 21797 => "1001010110001100", 21798 => "1111101000110010", 21799 => "1111011101101000", 21800 => "1001101001101110", 21801 => "1001010010110001", 21802 => "0111101011001011", 21803 => "0110011010001101", 21804 => "1100110010000001", 21805 => "1001010010100010", 21806 => "1001001010111110", 21807 => "1110101011011100", 21808 => "1000010111010100", 21809 => "1010110111010001", 21810 => "1111010000011101", 21811 => "0100000100100100", 21812 => "0101101000010111", 21813 => "0100101111110110", 21814 => "0011000110101000", 21815 => "0110110001101011", 21816 => "1110110100100010", 21817 => "1111110011111001", 21818 => "0010110111011001", 21819 => "1100101111001111", 21820 => "1111011101110110", 21821 => "1010001011000101", 21822 => "1110011101110101", 21823 => "1010100000101010", 21824 => "1011101101111101", 21825 => "1011101010000100", 21826 => "0010010001010100", 21827 => "1111011110001010", 21828 => "0011100010000011", 21829 => "1001011000101000", 21830 => "0110111011011011", 21831 => "0010001000001001", 21832 => "1110001011010111", 21833 => "1001011010111111", 21834 => "1101100000011100", 21835 => "0010111101011000", 21836 => "0101101011110110", 21837 => "0110001100001000", 21838 => "0000011000001001", 21839 => "1111100000110101", 21840 => "0100100001100011", 21841 => "1001010001111011", 21842 => "0111011101111001", 21843 => "0101101000010010", 21844 => "0010100010000010", 21845 => "1001011011111010", 21846 => "0010010000010111", 21847 => "1110010001101000", 21848 => "0110011111000100", 21849 => "1000100000111100", 21850 => "0110001001101111", 21851 => "0100000000010101", 21852 => "1110100011111110", 21853 => "0000000011100011", 21854 => "0111101011100110", 21855 => "0100010101010111", 21856 => "1010110101101111", 21857 => "0011010101001110", 21858 => "1111010111001001", 21859 => "0000011011110110", 21860 => "1110111000010011", 21861 => "1001100111111010", 21862 => "0001010011000011", 21863 => "1111110100101111", 21864 => "0111010011010000", 21865 => "0010011100001010", 21866 => "0100110101011110", 21867 => "1110101011010010", 21868 => "1101000100100000", 21869 => "1001000010110110", 21870 => "1111111101010110", 21871 => "0110111010000111", 21872 => "1000110101001001", 21873 => "0001101110010000", 21874 => "0001100111101011", 21875 => "0011100010110101", 21876 => "0010010001110111", 21877 => "1001101000010101", 21878 => "1001111010100000", 21879 => "1000100010110100", 21880 => "0110111000001111", 21881 => "0100101000101000", 21882 => "0001010000000100", 21883 => "1110011010101111", 21884 => "1001011010101111", 21885 => "0110010000011010", 21886 => "1010100110100000", 21887 => "1111000111100101", 21888 => "1101111100000010", 21889 => "0011001001001111", 21890 => "1001000110000100", 21891 => "0101110111110001", 21892 => "1100010011011100", 21893 => "1101001011110010", 21894 => "0101111101011000", 21895 => "1101010000111000", 21896 => "0100010111000100", 21897 => "1001110110010010", 21898 => "0000011000000100", 21899 => "0111001111010011", 21900 => "1010110011111011", 21901 => "0010110010000100", 21902 => "0001110011101001", 21903 => "0010001100100000", 21904 => "1101001111101010", 21905 => "1000010000101101", 21906 => "0111011000101110", 21907 => "1111001011010000", 21908 => "1001000110101101", 21909 => "1110110101110110", 21910 => "0110100001010010", 21911 => "0011010010100101", 21912 => "1001111101101110", 21913 => "1001000010000111", 21914 => "1100011001101111", 21915 => "0010010100101100", 21916 => "1011001100011000", 21917 => "1101110110011010", 21918 => "1100011010100010", 21919 => "1010111110100111", 21920 => "0000100101100111", 21921 => "0101110000101110", 21922 => "1111100110001000", 21923 => "1000001110011000", 21924 => "0001000011000000", 21925 => "1111010011000010", 21926 => "1111111111001011", 21927 => "0000010100101011", 21928 => "1010000110001011", 21929 => "1000111010101111", 21930 => "0110011101011000", 21931 => "0101100010101010", 21932 => "1110100111111010", 21933 => "0001111111100101", 21934 => "0100100101111110", 21935 => "0110100010011100", 21936 => "1110010101010100", 21937 => "0001011011110000", 21938 => "1111000101110000", 21939 => "0011000101100111", 21940 => "0111000000110010", 21941 => "0001001001010011", 21942 => "1101011110011000", 21943 => "0000010010000000", 21944 => "1110110010101001", 21945 => "1100011110101001", 21946 => "1101010010000101", 21947 => "1001000101111001", 21948 => "0011001010000001", 21949 => "0101111000010001", 21950 => "1101111100000000", 21951 => "1011011101101101", 21952 => "0011010011110000", 21953 => "0011111101100110", 21954 => "0101001011011101", 21955 => "0100010000010101", 21956 => "0011101101110001", 21957 => "0110110010001110", 21958 => "0100001000111010", 21959 => "1000000010011110", 21960 => "0001111101011000", 21961 => "1010100100101100", 21962 => "0110001011101011", 21963 => "1100000010101000", 21964 => "0011101001001101", 21965 => "0001101011101100", 21966 => "1110100001111110", 21967 => "0011111110011011", 21968 => "1001110100101000", 21969 => "1101110011111001", 21970 => "1100001111011001", 21971 => "0011010100100101", 21972 => "1111011111101011", 21973 => "1011110011010101", 21974 => "0110110110110100", 21975 => "0110010100010010", 21976 => "0001100010001000", 21977 => "1011010111100000", 21978 => "0001000001011001", 21979 => "0000010000010000", 21980 => "0101110111100010", 21981 => "0110001001101000", 21982 => "0110001010101100", 21983 => "1011111001100000", 21984 => "1111101110101110", 21985 => "0011010111111111", 21986 => "0001101100001010", 21987 => "1010011111010011", 21988 => "0001110011100000", 21989 => "0100111000010001", 21990 => "1000001110100010", 21991 => "1001110100111100", 21992 => "1011010011011100", 21993 => "0011100101101111", 21994 => "0011100000111111", 21995 => "1001100011100100", 21996 => "1011110010100110", 21997 => "1100000001100010", 21998 => "1100000101100101", 21999 => "0110100110010101", 22000 => "0101001011110001", 22001 => "0101100101011111", 22002 => "0000000011110001", 22003 => "0101010000010001", 22004 => "1011101110010011", 22005 => "1010110011001000", 22006 => "1111101111111110", 22007 => "0010001010111011", 22008 => "1110011011011100", 22009 => "0010001000100111", 22010 => "1000011101011010", 22011 => "0010011110010111", 22012 => "1100111111110101", 22013 => "1101111100000001", 22014 => "0010010100011011", 22015 => "0111000011101100", 22016 => "0100100001100011", 22017 => "1010000101011000", 22018 => "1010111101110101", 22019 => "0101111110011010", 22020 => "0011011100110101", 22021 => "0100111000100111", 22022 => "0011010110001110", 22023 => "0001001001111010", 22024 => "0000001101111110", 22025 => "0111001010000011", 22026 => "1110000101100101", 22027 => "1100001100000010", 22028 => "1101101101101001", 22029 => "0110010000010101", 22030 => "1011000010101010", 22031 => "1101110011000011", 22032 => "0100100100001001", 22033 => "1101001100000110", 22034 => "0001101111000101", 22035 => "0010100011100011", 22036 => "0001101110000111", 22037 => "0001010001111010", 22038 => "1000100100001110", 22039 => "0100011001111011", 22040 => "1101000101000011", 22041 => "0110000011110100", 22042 => "0110010000001010", 22043 => "1101101110001010", 22044 => "0001110100010111", 22045 => "0001010110100110", 22046 => "0011001001010101", 22047 => "1101001101000001", 22048 => "1011000000000101", 22049 => "0100010011010111", 22050 => "1111101001001101", 22051 => "1101101111001110", 22052 => "1001010100110100", 22053 => "0000011010010101", 22054 => "1101100100001000", 22055 => "0001110010111001", 22056 => "0011110001000111", 22057 => "1101011100110011", 22058 => "0101110100000011", 22059 => "0011001110010100", 22060 => "0110001000100000", 22061 => "1101100001110010", 22062 => "0111100011111001", 22063 => "0111110110010111", 22064 => "0101110010001001", 22065 => "0100000011101111", 22066 => "1100000111001100", 22067 => "1110000111101111", 22068 => "1100100010101001", 22069 => "1100100101111001", 22070 => "1011000100000011", 22071 => "0100001011001000", 22072 => "0011010111001110", 22073 => "1101011001001111", 22074 => "1101101011011011", 22075 => "0000101101111001", 22076 => "1010111001111010", 22077 => "1011001000101010", 22078 => "1111001111111001", 22079 => "0110101110100110", 22080 => "0001101001110010", 22081 => "1010000110110101", 22082 => "1110001100010011", 22083 => "1000001110110110", 22084 => "0101110011110111", 22085 => "1010111011111001", 22086 => "1100010111010011", 22087 => "0101100110111000", 22088 => "0111110110111110", 22089 => "0101110100010011", 22090 => "1000011101100001", 22091 => "1001101001001010", 22092 => "1001110111100101", 22093 => "1100100101010100", 22094 => "0010011001101001", 22095 => "0000101110001110", 22096 => "1001010000111011", 22097 => "1100000010111111", 22098 => "0011111111000000", 22099 => "0110110011001010", 22100 => "1100110110111111", 22101 => "0000010101000110", 22102 => "1100011101001011", 22103 => "1010001101010010", 22104 => "1100111111011111", 22105 => "1100111111101110", 22106 => "0100000100111100", 22107 => "0001000001100111", 22108 => "0011011010101100", 22109 => "1100110001000000", 22110 => "0111011000010001", 22111 => "1111011011011010", 22112 => "0110111011011110", 22113 => "1001111101010011", 22114 => "1110010001000000", 22115 => "0110011000010001", 22116 => "1001010100010100", 22117 => "1111100111010000", 22118 => "0100000111000010", 22119 => "0011110111001101", 22120 => "1111101100111100", 22121 => "1111101110110000", 22122 => "0011100000110010", 22123 => "1000110111111101", 22124 => "0101000001111011", 22125 => "1000111100100100", 22126 => "1011001001001010", 22127 => "1001100000101001", 22128 => "1100110000000001", 22129 => "0101110010011111", 22130 => "1110100010011101", 22131 => "1111100100110100", 22132 => "0110111010000100", 22133 => "1111101101011110", 22134 => "0011101010000101", 22135 => "1111110110010011", 22136 => "1101001111100110", 22137 => "0011011011010011", 22138 => "0000010111110000", 22139 => "0100100010001101", 22140 => "1011001101101011", 22141 => "1001111111001111", 22142 => "1011011011010011", 22143 => "0010001010110011", 22144 => "1100100100010000", 22145 => "0011001110001010", 22146 => "0111111010010010", 22147 => "0011011100111011", 22148 => "1111100011111100", 22149 => "1011011101111100", 22150 => "0001010110100111", 22151 => "0101001110010100", 22152 => "0011011000100110", 22153 => "0111001111000000", 22154 => "1001011000011101", 22155 => "0010110011110100", 22156 => "0101010110100110", 22157 => "0001001001000110", 22158 => "0000000100101111", 22159 => "1010001101000001", 22160 => "0110011110000110", 22161 => "1100101001110011", 22162 => "1001111110010011", 22163 => "1110100111111010", 22164 => "0010001110111111", 22165 => "0110110011110001", 22166 => "1111000101111011", 22167 => "0100010100010011", 22168 => "1101010011011110", 22169 => "0111011011110001", 22170 => "0111111000101000", 22171 => "0011001011001101", 22172 => "1001011010111000", 22173 => "1010111011100111", 22174 => "1011010111101101", 22175 => "1101110001011000", 22176 => "0101010000011110", 22177 => "1111000000010000", 22178 => "1101011011111000", 22179 => "0001100110011100", 22180 => "0000111111011100", 22181 => "1101111100111001", 22182 => "0010110000100000", 22183 => "1001100010110110", 22184 => "0000001100111001", 22185 => "1011101011000110", 22186 => "1100000100110000", 22187 => "0011000011010111", 22188 => "1111111110000011", 22189 => "0100001000011000", 22190 => "1000100010111000", 22191 => "0101001110100010", 22192 => "1100101001001011", 22193 => "0000011111100001", 22194 => "0110110110111100", 22195 => "0011101011100111", 22196 => "1111011101110110", 22197 => "0110111000000110", 22198 => "0100110010011111", 22199 => "0110000101001111", 22200 => "0101100000111100", 22201 => "1010001110000001", 22202 => "0110100011010101", 22203 => "1000110011111101", 22204 => "1010001000100010", 22205 => "0110011011100001", 22206 => "1111011010001111", 22207 => "1111010001011111", 22208 => "1111011010110110", 22209 => "1000001100110111", 22210 => "1011011011100011", 22211 => "1101101111011100", 22212 => "0000111100110000", 22213 => "1001111010110111", 22214 => "1011001110000100", 22215 => "1010001111100100", 22216 => "0011111110110011", 22217 => "0110100011101001", 22218 => "0111100000111110", 22219 => "0000101000000101", 22220 => "0101100000000001", 22221 => "1011000100100110", 22222 => "0010000010110100", 22223 => "0001100011001100", 22224 => "0001000111111001", 22225 => "0001011000010010", 22226 => "0100100100011000", 22227 => "1010100001101010", 22228 => "1000110011011100", 22229 => "1111110000000101", 22230 => "0110000111110100", 22231 => "0100111111010011", 22232 => "1100101011100111", 22233 => "1111110111001100", 22234 => "1100101010110100", 22235 => "1111001101100010", 22236 => "1110001101110000", 22237 => "1001001111100011", 22238 => "1010010001101100", 22239 => "0011101111111010", 22240 => "1101100010001110", 22241 => "1001100011100110", 22242 => "0010110100010100", 22243 => "0101110001110111", 22244 => "1110000100011101", 22245 => "1101000110100110", 22246 => "1010111101100111", 22247 => "0101001011100111", 22248 => "0011101110100001", 22249 => "0101001001001110", 22250 => "0000001000000100", 22251 => "0110000101111011", 22252 => "0110001000001110", 22253 => "0100000110111001", 22254 => "0111011111101001", 22255 => "1001000000111001", 22256 => "0101010101111001", 22257 => "1100000111001011", 22258 => "1010000101100010", 22259 => "0101001011111100", 22260 => "0001010011010111", 22261 => "0001111101100101", 22262 => "0010111011101110", 22263 => "1100111111000010", 22264 => "0110111100001000", 22265 => "1010010001111001", 22266 => "0111111010011101", 22267 => "0111110010111100", 22268 => "0010111011000100", 22269 => "1001110010101110", 22270 => "0011010100100110", 22271 => "0110101011001100", 22272 => "1001110100110001", 22273 => "0010101001111000", 22274 => "1001110100100000", 22275 => "0001110111010011", 22276 => "0111101000111001", 22277 => "1101100100101010", 22278 => "1010111000000101", 22279 => "1110100110101101", 22280 => "0001000101001011", 22281 => "0100010100111100", 22282 => "0100100011111100", 22283 => "0011101000110010", 22284 => "1000110010010111", 22285 => "0100101101101010", 22286 => "0001011111010000", 22287 => "0110000000000110", 22288 => "0101010000010000", 22289 => "0111110101101101", 22290 => "0001000010110101", 22291 => "1100110001001110", 22292 => "0100000000100001", 22293 => "0010001010101010", 22294 => "1000010101101110", 22295 => "0011010111100110", 22296 => "1100101001110010", 22297 => "0000001100111111", 22298 => "1101010110111111", 22299 => "1010110010011110", 22300 => "0011111101001001", 22301 => "0111001010001101", 22302 => "1001101001110000", 22303 => "1101100011101110", 22304 => "1111011100110011", 22305 => "0101111111010010", 22306 => "1100101000111101", 22307 => "1011010000111110", 22308 => "0100011000000001", 22309 => "1001011001011100", 22310 => "1110000111100001", 22311 => "0001011101000000", 22312 => "1101111101111000", 22313 => "1110100101100111", 22314 => "1011001110101010", 22315 => "0010000111000100", 22316 => "0010110101010000", 22317 => "1100100100001110", 22318 => "0111011110011101", 22319 => "0100111010111011", 22320 => "0101101101110001", 22321 => "0010011010100000", 22322 => "0010000100010110", 22323 => "0110010001011100", 22324 => "0011111010001100", 22325 => "0101011100101010", 22326 => "1100111010111011", 22327 => "1000110100101101", 22328 => "0101111010111001", 22329 => "0101110110101010", 22330 => "1110010001000110", 22331 => "0111000010000101", 22332 => "0000101001011101", 22333 => "0001111001011011", 22334 => "0100110100010111", 22335 => "1001110010000000", 22336 => "1001101010110111", 22337 => "1110111010111111", 22338 => "1001001010111111", 22339 => "1010010101010011", 22340 => "1001101111100001", 22341 => "0100111110011000", 22342 => "1110100000000110", 22343 => "0001010010110001", 22344 => "0011101000111010", 22345 => "1011100101100110", 22346 => "1101000101111001", 22347 => "0011101011110010", 22348 => "0110100100000010", 22349 => "1100011010111110", 22350 => "1001110011110000", 22351 => "0100101100001110", 22352 => "0001011101101110", 22353 => "1111100010000110", 22354 => "1101101111001011", 22355 => "1110111000011111", 22356 => "0001110110101100", 22357 => "1100100011000011", 22358 => "0010110011011111", 22359 => "1011010010010011", 22360 => "1110111011011001", 22361 => "1010100100001001", 22362 => "1000110010110110", 22363 => "0011001010110011", 22364 => "1100001011111100", 22365 => "1110100100100111", 22366 => "1111000111001111", 22367 => "1110100101101000", 22368 => "1100011000101011", 22369 => "1011101001110011", 22370 => "0011001010010010", 22371 => "0001001101100101", 22372 => "1101101110011101", 22373 => "0011101100100010", 22374 => "1111100101110100", 22375 => "0110001101101100", 22376 => "0111001011111000", 22377 => "1000110011111110", 22378 => "0000010001110000", 22379 => "0100011001010110", 22380 => "0010001111011000", 22381 => "0100110111010010", 22382 => "1000101010100011", 22383 => "1000010001110100", 22384 => "0101110101111000", 22385 => "1101100101100010", 22386 => "1111010111000110", 22387 => "0011110101010101", 22388 => "0011010111010011", 22389 => "1001010010001110", 22390 => "1000111110110001", 22391 => "0101011011000110", 22392 => "0101010110100001", 22393 => "0111100111011110", 22394 => "1001101111111101", 22395 => "0011101110110001", 22396 => "1100111101010001", 22397 => "0010010110110110", 22398 => "1111010110001001", 22399 => "1111011000010111", 22400 => "1101000010001101", 22401 => "1100000010001011", 22402 => "1111011010010110", 22403 => "1101011001110100", 22404 => "1110110111000101", 22405 => "0001000100000010", 22406 => "0001110110001001", 22407 => "1010100000111011", 22408 => "1110011011111000", 22409 => "0000001001111111", 22410 => "1101110100110111", 22411 => "1000010001000101", 22412 => "1101001101000101", 22413 => "0101110011110101", 22414 => "0011011010110111", 22415 => "0001111110011000", 22416 => "1111110011100111", 22417 => "0100011110010010", 22418 => "1100100000011101", 22419 => "0100101101101100", 22420 => "1011001111111011", 22421 => "0101101001111011", 22422 => "0101011000010111", 22423 => "0001111110000111", 22424 => "1110001110101010", 22425 => "1000101101100111", 22426 => "0000010001110101", 22427 => "1011001001010011", 22428 => "0100011110000100", 22429 => "0001100100000010", 22430 => "0101101001001010", 22431 => "0100011100100100", 22432 => "1100010111111100", 22433 => "1110111000101100", 22434 => "1110101110111111", 22435 => "1000101100010100", 22436 => "0001000111110110", 22437 => "1010011100000010", 22438 => "0110100110101000", 22439 => "0101000011111100", 22440 => "0111111111001011", 22441 => "0000111110101001", 22442 => "1111101111000100", 22443 => "1111011001100000", 22444 => "1111000001111000", 22445 => "0000000110101100", 22446 => "1100110100110101", 22447 => "1010010001111111", 22448 => "0111010011100100", 22449 => "1001010101100111", 22450 => "1011101010000001", 22451 => "1101110000010011", 22452 => "0001101011101101", 22453 => "1100101010111111", 22454 => "0110101000110100", 22455 => "0000011100101000", 22456 => "1100011001110101", 22457 => "0100001010101011", 22458 => "1010001011100000", 22459 => "1100100110111011", 22460 => "0111010101010000", 22461 => "0001011110100101", 22462 => "0100101001111000", 22463 => "0001011010001111", 22464 => "1011101011000110", 22465 => "1000110000000011", 22466 => "1110010100111100", 22467 => "0010001001111001", 22468 => "1111001001010000", 22469 => "0011101101001110", 22470 => "1001011101110100", 22471 => "1000111011011110", 22472 => "0000101100110001", 22473 => "1010010011000101", 22474 => "1100010111011011", 22475 => "0101010001101000", 22476 => "1000001010111000", 22477 => "0000011101001000", 22478 => "0111010010000001", 22479 => "1111101011110011", 22480 => "0101101010010000", 22481 => "0000010001110101", 22482 => "1110001101110110", 22483 => "0111000001111101", 22484 => "1000001111011110", 22485 => "0110100010110100", 22486 => "0111001101111110", 22487 => "1010111100101110", 22488 => "1101110001111000", 22489 => "0000010110101111", 22490 => "1100001100100011", 22491 => "0101011110101110", 22492 => "1000101111010011", 22493 => "0001100010111000", 22494 => "0101010011100001", 22495 => "1110100101011101", 22496 => "1001111111000111", 22497 => "1011111001101111", 22498 => "1000100011111111", 22499 => "0110011101111000", 22500 => "0110001000111100", 22501 => "1001100000010111", 22502 => "0111001100111101", 22503 => "1011101000000001", 22504 => "1101001010001011", 22505 => "0101100010110101", 22506 => "1001110111111000", 22507 => "1001111000111111", 22508 => "0100011000001010", 22509 => "0011100001001010", 22510 => "1000110001000100", 22511 => "1000101111110101", 22512 => "1110010010000101", 22513 => "0010010111110010", 22514 => "1010111001000110", 22515 => "1101110001001000", 22516 => "0100100110101111", 22517 => "0000101010010000", 22518 => "1100010100100001", 22519 => "1111011000111001", 22520 => "1011111100010011", 22521 => "1100110011011010", 22522 => "0011110110100111", 22523 => "0010100110011100", 22524 => "0011100010001010", 22525 => "1100011101111111", 22526 => "0101111010111101", 22527 => "0011011100001100", 22528 => "0000011010110110", 22529 => "1010010001110111", 22530 => "0010101110010110", 22531 => "0101111011111110", 22532 => "0110100000001010", 22533 => "0101111100010010", 22534 => "0101011001011111", 22535 => "1110010001111101", 22536 => "0010000111000111", 22537 => "0010000000000011", 22538 => "1100110100110000", 22539 => "0000001111110100", 22540 => "0001101100010011", 22541 => "1000100001100001", 22542 => "0111110100001000", 22543 => "0010000100100000", 22544 => "1101100011110000", 22545 => "1100001001011001", 22546 => "0000001111011011", 22547 => "0010010100001111", 22548 => "0110111101100011", 22549 => "0001101011100100", 22550 => "0011101110111000", 22551 => "0111000101100101", 22552 => "0101000111110100", 22553 => "1001000101011100", 22554 => "1011110000010111", 22555 => "1001100001101010", 22556 => "0000100111010000", 22557 => "0010011001010001", 22558 => "1100000110011110", 22559 => "0111100101011110", 22560 => "0111010110010111", 22561 => "0110000100110001", 22562 => "1111011111011110", 22563 => "1100000011001011", 22564 => "1100000011010110", 22565 => "0000110111101001", 22566 => "1010111111100111", 22567 => "1010011001101110", 22568 => "0101111100011111", 22569 => "1011110110101000", 22570 => "0010100000000101", 22571 => "0000010100000010", 22572 => "1010000110011011", 22573 => "1111111110111100", 22574 => "0101100011000110", 22575 => "0001010001111101", 22576 => "1101110110111101", 22577 => "1000101011101110", 22578 => "0100101011110110", 22579 => "1001110111101001", 22580 => "0100110010100010", 22581 => "1110011010000111", 22582 => "0000010111011000", 22583 => "0110000100000110", 22584 => "0101111010011100", 22585 => "0110011110010100", 22586 => "0011001000010110", 22587 => "1101000111110110", 22588 => "0100001000000010", 22589 => "1001011010010010", 22590 => "0011101100011000", 22591 => "1110100011111100", 22592 => "1101110011010111", 22593 => "0110001011001011", 22594 => "1110001000111100", 22595 => "1100001011100101", 22596 => "1110011010001110", 22597 => "1101001010100000", 22598 => "0100100101001011", 22599 => "1011001011001000", 22600 => "0011101101111000", 22601 => "0100111010000010", 22602 => "0001100111011100", 22603 => "1101010100011011", 22604 => "0011100001000101", 22605 => "0000100001100001", 22606 => "0100100101101000", 22607 => "1001110100000011", 22608 => "0111100000101111", 22609 => "1000001010010110", 22610 => "1000100010001110", 22611 => "1110100000001001", 22612 => "1100101111010001", 22613 => "0100010001010110", 22614 => "0110001111101011", 22615 => "0010111011111111", 22616 => "1110100000101011", 22617 => "1111111101001110", 22618 => "0000100100011111", 22619 => "1011001011111100", 22620 => "1011110100001110", 22621 => "1001110010100011", 22622 => "0000101110101001", 22623 => "1000011111011111", 22624 => "1111001101000010", 22625 => "0101101100011111", 22626 => "1001001011001100", 22627 => "0110001110000101", 22628 => "1011010001000000", 22629 => "1100000000000001", 22630 => "1001000000000111", 22631 => "0000110000111111", 22632 => "1101010000010011", 22633 => "0011010001111111", 22634 => "0011010001101110", 22635 => "0001100110011000", 22636 => "0101110000111010", 22637 => "1010000001110011", 22638 => "0110001010001110", 22639 => "0010110101001001", 22640 => "0111100011101111", 22641 => "1100010001000010", 22642 => "1000101111011110", 22643 => "0010111000111010", 22644 => "0111111111000001", 22645 => "0011000110000100", 22646 => "1101010101001101", 22647 => "1011101111100111", 22648 => "0110001110110011", 22649 => "1111110101110000", 22650 => "0100111111111001", 22651 => "1110111101011100", 22652 => "0100011000111101", 22653 => "1101000011100111", 22654 => "0001000111100110", 22655 => "0110000000101100", 22656 => "0010011010110000", 22657 => "0110001101010111", 22658 => "1110100101010111", 22659 => "1110001101100111", 22660 => "1110001000010001", 22661 => "1010010000001000", 22662 => "1001010001000010", 22663 => "1011101000111101", 22664 => "0100101110100011", 22665 => "0000110100110010", 22666 => "0010001011010101", 22667 => "1001110111011000", 22668 => "1111001010010001", 22669 => "1110010100100100", 22670 => "1010110000101110", 22671 => "1100111011100100", 22672 => "0011011111111101", 22673 => "0110001000000000", 22674 => "0000011000111000", 22675 => "0101101001110001", 22676 => "1100010000110111", 22677 => "1010100011111011", 22678 => "0001001001111001", 22679 => "1111000110001111", 22680 => "0000001100101000", 22681 => "0110100000001000", 22682 => "1100000010011000", 22683 => "0100001101011111", 22684 => "0101000001001110", 22685 => "1000010111110011", 22686 => "1010100000111010", 22687 => "0100010111101101", 22688 => "0010110101011101", 22689 => "1010000000010010", 22690 => "0111101001011100", 22691 => "0111111100010000", 22692 => "0001100000100100", 22693 => "1001110100001001", 22694 => "0000011111000000", 22695 => "1100001011001001", 22696 => "0110101101100101", 22697 => "0011100100100111", 22698 => "1100010111011001", 22699 => "0100000111011010", 22700 => "1011101010111101", 22701 => "1101010110000000", 22702 => "1100011010001011", 22703 => "0000110010100010", 22704 => "1100101110010110", 22705 => "0001101001010001", 22706 => "0101000100010101", 22707 => "0100111001111011", 22708 => "0101111101010010", 22709 => "0111001100000100", 22710 => "0111001010011000", 22711 => "1000111001001001", 22712 => "1110101011010011", 22713 => "1101101110101110", 22714 => "0000001000111001", 22715 => "0011101101111101", 22716 => "0001100000100100", 22717 => "1011000101000000", 22718 => "1000100000111110", 22719 => "0110110010110110", 22720 => "1000101010110101", 22721 => "1001101001011111", 22722 => "0110100010110101", 22723 => "0110101010110100", 22724 => "1111000110011110", 22725 => "0001111100001111", 22726 => "1000100010011111", 22727 => "0111101100100000", 22728 => "0011100011100100", 22729 => "0100110011110010", 22730 => "0111110100110100", 22731 => "0100000010111001", 22732 => "1111110111100110", 22733 => "0001110000000000", 22734 => "0101100001101100", 22735 => "1001111011000101", 22736 => "1101111010101101", 22737 => "0101000110001010", 22738 => "0111011100010110", 22739 => "1011110000110100", 22740 => "1111010001110000", 22741 => "0011110000101010", 22742 => "0001001001100001", 22743 => "1111001001000111", 22744 => "0010111001011011", 22745 => "1011111011101010", 22746 => "0011111111110101", 22747 => "0101011011110000", 22748 => "1001011101001011", 22749 => "1001111011011001", 22750 => "1001010111100001", 22751 => "0001100101010101", 22752 => "1000100100010101", 22753 => "0100010110001001", 22754 => "0010110101111001", 22755 => "0111001000101001", 22756 => "1010111100111100", 22757 => "1010011001101110", 22758 => "1011100111110010", 22759 => "0010111100111001", 22760 => "0110111110100110", 22761 => "0110100101000010", 22762 => "1001101101111010", 22763 => "0110100110100101", 22764 => "1011101010011111", 22765 => "1100010011011010", 22766 => "0000100010111101", 22767 => "0100001101011000", 22768 => "0001111010001101", 22769 => "0110011001001101", 22770 => "0110011110110100", 22771 => "1010011110010110", 22772 => "0111101010010101", 22773 => "1111110011101101", 22774 => "0011101000000011", 22775 => "1000110010011010", 22776 => "0010011010010001", 22777 => "1100110011011111", 22778 => "0011011110110001", 22779 => "0110010000110101", 22780 => "1000100110000001", 22781 => "0000100010100111", 22782 => "0111100001100110", 22783 => "0111011011011111", 22784 => "1010001110011000", 22785 => "1001100001000101", 22786 => "1011010011111011", 22787 => "0111010011101001", 22788 => "0100000111111111", 22789 => "1111100010001100", 22790 => "0110111111000000", 22791 => "1000010101000100", 22792 => "0100011000010110", 22793 => "1001010111001101", 22794 => "0111101011001100", 22795 => "1000010100110110", 22796 => "1101100111110010", 22797 => "1011110011010101", 22798 => "1000010110011101", 22799 => "1110001010001100", 22800 => "0001001010111000", 22801 => "1010100110110001", 22802 => "1110100001110010", 22803 => "0101001001100101", 22804 => "0010011110111010", 22805 => "1011101101110110", 22806 => "0111111000000100", 22807 => "0100100110010111", 22808 => "0111001000011011", 22809 => "1101111100001100", 22810 => "0011010001000110", 22811 => "1110111101101110", 22812 => "1001000100111011", 22813 => "1100000000011100", 22814 => "1000011111010000", 22815 => "0011100010011000", 22816 => "0001000110001110", 22817 => "1111010110100100", 22818 => "1100100101011111", 22819 => "1000011000101000", 22820 => "1100011000011011", 22821 => "0000101101011110", 22822 => "1011110100111001", 22823 => "1011111001100010", 22824 => "1100101111110100", 22825 => "0011101001101111", 22826 => "1110010011011000", 22827 => "1001001010010100", 22828 => "0101000010111000", 22829 => "1101110110110101", 22830 => "1000111010100110", 22831 => "1111100100100011", 22832 => "0011011011010010", 22833 => "1100101010011100", 22834 => "0100111100111001", 22835 => "1001010001101110", 22836 => "1011101010010010", 22837 => "0001110110001110", 22838 => "1111001100010000", 22839 => "1110001000010001", 22840 => "0011010000101011", 22841 => "0100101000000101", 22842 => "0010110000011111", 22843 => "1011011111000110", 22844 => "1111110101111100", 22845 => "1011100001101111", 22846 => "0111001110001110", 22847 => "0001001011111100", 22848 => "0110011011100011", 22849 => "1000000000001000", 22850 => "1010000100011001", 22851 => "0001001111110001", 22852 => "0010111011010101", 22853 => "1010000011101010", 22854 => "1111011111110111", 22855 => "1010110000100011", 22856 => "0101110110000101", 22857 => "0011110101111101", 22858 => "0111111101110110", 22859 => "0011010110000001", 22860 => "0110110000011010", 22861 => "1001000110111011", 22862 => "1111010101101011", 22863 => "1110001100100010", 22864 => "0001010000100100", 22865 => "1000110100000110", 22866 => "1100011111111001", 22867 => "1000000010100000", 22868 => "0111001000011000", 22869 => "1001110101001000", 22870 => "0000101011011111", 22871 => "0001101000011100", 22872 => "0110111001011111", 22873 => "1111111101110110", 22874 => "1100111001011110", 22875 => "0011011111100010", 22876 => "1011000000110100", 22877 => "0010100000010110", 22878 => "0000100100011001", 22879 => "0111101011111111", 22880 => "0010101000000010", 22881 => "1000101110011100", 22882 => "1010101000101000", 22883 => "1111111110111000", 22884 => "0000110010100101", 22885 => "1001110000001000", 22886 => "0100010001100111", 22887 => "1111100100010101", 22888 => "1011100110000001", 22889 => "1100001111110111", 22890 => "1000101111110011", 22891 => "1010111000111111", 22892 => "1000011011101111", 22893 => "1100110101010111", 22894 => "1001010011011001", 22895 => "0010100111010000", 22896 => "0101101111110001", 22897 => "1110111110011100", 22898 => "1111001110011100", 22899 => "0101001011011110", 22900 => "0111100010000101", 22901 => "0101001101101010", 22902 => "1010100001100011", 22903 => "1110111100100001", 22904 => "0100111000010001", 22905 => "1001110110111011", 22906 => "1001110010101001", 22907 => "0000010110100111", 22908 => "1101010000101101", 22909 => "0101010010001011", 22910 => "1110010100110111", 22911 => "0111001100000001", 22912 => "0000101100111101", 22913 => "1111100001010001", 22914 => "0000101101111010", 22915 => "0101010110000000", 22916 => "1000010000100000", 22917 => "1101001110100101", 22918 => "1100000010101000", 22919 => "1111101100101001", 22920 => "0110001011001001", 22921 => "0111100101110000", 22922 => "0001100101000001", 22923 => "1110101010101001", 22924 => "0101110100100100", 22925 => "1111000110011011", 22926 => "1001111100000100", 22927 => "1100010011101000", 22928 => "0011100101000000", 22929 => "1110100111000010", 22930 => "1001000010000110", 22931 => "0110000000010010", 22932 => "1101111101110101", 22933 => "1000101010001110", 22934 => "0001110111101010", 22935 => "0100010011001010", 22936 => "0001001101001000", 22937 => "1110011000101100", 22938 => "0100001101011011", 22939 => "1110101010011000", 22940 => "0001000101001111", 22941 => "1001111001111000", 22942 => "1110100101001101", 22943 => "0101001000100010", 22944 => "1001000000111001", 22945 => "1000110111011100", 22946 => "1001000110110100", 22947 => "0001100011011100", 22948 => "0100101011011011", 22949 => "0110010000100011", 22950 => "0011010100110011", 22951 => "0100011001110010", 22952 => "1011101100101011", 22953 => "0010000010100100", 22954 => "0111011101001000", 22955 => "1010110101011010", 22956 => "1110101001110110", 22957 => "0000001001110111", 22958 => "0011011000011010", 22959 => "1111101000001101", 22960 => "1000101110001001", 22961 => "0000000010110110", 22962 => "1001110100110001", 22963 => "1101010001100100", 22964 => "0111111111010101", 22965 => "1011101001000011", 22966 => "0010000100010001", 22967 => "0101110000010110", 22968 => "1110001001001001", 22969 => "0010010101010010", 22970 => "0001000100110111", 22971 => "0101100100000010", 22972 => "0000111010011011", 22973 => "1101000110001001", 22974 => "0001010110101101", 22975 => "0001011001000111", 22976 => "1100001000101100", 22977 => "0101101000010001", 22978 => "0011101000000111", 22979 => "0011011011111000", 22980 => "1101110111001000", 22981 => "1101011000110100", 22982 => "1010001010100001", 22983 => "1101110001110111", 22984 => "1000001001101110", 22985 => "0100010100111000", 22986 => "1101110111011010", 22987 => "0111001100101001", 22988 => "1101100010010110", 22989 => "1101011101001011", 22990 => "1000100100100010", 22991 => "0100100010111111", 22992 => "0010001101010001", 22993 => "1101011011011101", 22994 => "0111011111000001", 22995 => "1001101001111011", 22996 => "1001101101000100", 22997 => "0100011000110111", 22998 => "0110001010001100", 22999 => "0100001010000010", 23000 => "1001011101110010", 23001 => "1001100100111100", 23002 => "1101001000000000", 23003 => "1000001100100111", 23004 => "1000100001110010", 23005 => "0110000100100010", 23006 => "1100010000000101", 23007 => "1111001011011111", 23008 => "0101100111111110", 23009 => "0111111111010010", 23010 => "1110101101010010", 23011 => "1000000010101010", 23012 => "1110111101101000", 23013 => "1001001000010010", 23014 => "0010101011110111", 23015 => "0110101101000011", 23016 => "0100101000010111", 23017 => "1111000000110100", 23018 => "0001001011011111", 23019 => "0111111101001110", 23020 => "0101111111001101", 23021 => "0111100101001100", 23022 => "0111111110000010", 23023 => "0100011111011100", 23024 => "1101001000101010", 23025 => "1100101000001111", 23026 => "0001100100101001", 23027 => "1001101000101100", 23028 => "1100001110010000", 23029 => "0001001011111110", 23030 => "0101100011011000", 23031 => "1001111110000001", 23032 => "0110110111010001", 23033 => "0000001011110011", 23034 => "1001101101111000", 23035 => "1110110111111111", 23036 => "0100010000100110", 23037 => "0001010011000101", 23038 => "1010011111111100", 23039 => "1010011111010000", 23040 => "1010101000010000", 23041 => "1010100110110000", 23042 => "1000001101101010", 23043 => "1111011111011100", 23044 => "0010011001101111", 23045 => "1101110110001111", 23046 => "1001001101000000", 23047 => "1010111110011001", 23048 => "1100111000100000", 23049 => "0100100111010101", 23050 => "1111000111101110", 23051 => "1010001101011011", 23052 => "1101110011010111", 23053 => "1100010000100010", 23054 => "0010111101100010", 23055 => "0000010110111010", 23056 => "0101011010101111", 23057 => "1011011100000111", 23058 => "1001101110101000", 23059 => "1100001001010101", 23060 => "1000000110111010", 23061 => "0001100010101011", 23062 => "0001000100110111", 23063 => "0001010100001100", 23064 => "0111001011111101", 23065 => "1010100101101011", 23066 => "1001010111111011", 23067 => "0110111111001011", 23068 => "0110011000110100", 23069 => "1101001000111010", 23070 => "0111011000001001", 23071 => "0000111000100001", 23072 => "0101000010110000", 23073 => "1100011100100101", 23074 => "0111010000100010", 23075 => "0101100000101011", 23076 => "1100110010011001", 23077 => "0111000110000001", 23078 => "1010101000100110", 23079 => "1100011101111000", 23080 => "1100010000001000", 23081 => "1110001010111111", 23082 => "0001111111111010", 23083 => "0000011011100110", 23084 => "0100110011100101", 23085 => "1000100000010100", 23086 => "1000111001000100", 23087 => "0110001100000100", 23088 => "0010110000110101", 23089 => "1101001110001111", 23090 => "1000100010010011", 23091 => "1100111100111101", 23092 => "0111101101001101", 23093 => "0010000001100010", 23094 => "0001001100011010", 23095 => "0110100000011001", 23096 => "0110001110000010", 23097 => "0110100111000000", 23098 => "1010111011111000", 23099 => "1101011100101000", 23100 => "0110010101111111", 23101 => "1011101110011101", 23102 => "0101000100010000", 23103 => "1010001001110011", 23104 => "0011001111101001", 23105 => "0000000000000110", 23106 => "0100100001110110", 23107 => "1000110100000100", 23108 => "0010101010110000", 23109 => "0111001010111000", 23110 => "1101100110100001", 23111 => "1011001100101001", 23112 => "0110000011011101", 23113 => "0101011101110111", 23114 => "1111010101000101", 23115 => "1011110000000001", 23116 => "1010011111111010", 23117 => "0100010000001011", 23118 => "0001000100110101", 23119 => "1011101000100010", 23120 => "1010110110101111", 23121 => "0001001011100011", 23122 => "0101110101100001", 23123 => "0101101111101000", 23124 => "0000111111110001", 23125 => "0111000111000001", 23126 => "0101000010001000", 23127 => "0100110010110101", 23128 => "0011010101001001", 23129 => "1001100001100111", 23130 => "0000010001000001", 23131 => "0000010011001010", 23132 => "1001110110100011", 23133 => "0101110100100111", 23134 => "1101111010010111", 23135 => "0000111100111001", 23136 => "1100000010000010", 23137 => "0101000101010011", 23138 => "0010000011101100", 23139 => "0001001111110011", 23140 => "1110011100111000", 23141 => "0100000111111010", 23142 => "1011100011001001", 23143 => "0011111110010000", 23144 => "1111010010010010", 23145 => "0100110010111111", 23146 => "0000111111111110", 23147 => "1001000110010011", 23148 => "1101101110010111", 23149 => "0001000111101000", 23150 => "0010000001101101", 23151 => "0001110001001101", 23152 => "0010101000001111", 23153 => "1100000010111001", 23154 => "1101110100001010", 23155 => "0000011110100110", 23156 => "1000100000100111", 23157 => "0011111110000010", 23158 => "0101110111001101", 23159 => "0010010000111001", 23160 => "0011000000000001", 23161 => "1000000000110010", 23162 => "1011011011100111", 23163 => "1110111110110111", 23164 => "0010000000111100", 23165 => "1100000000110011", 23166 => "1000111011000010", 23167 => "0000011110111100", 23168 => "0101011100111001", 23169 => "0101110001010010", 23170 => "0000110111001010", 23171 => "1111010110110001", 23172 => "0011001001010101", 23173 => "1100110111111100", 23174 => "1110010100110010", 23175 => "0100110010000101", 23176 => "1111010100100000", 23177 => "0000010100111110", 23178 => "0111101100101111", 23179 => "0001111110010110", 23180 => "0111001100010100", 23181 => "1010001101110111", 23182 => "0000010011010111", 23183 => "0110010110110111", 23184 => "0011101010101100", 23185 => "1100101110011111", 23186 => "0110011101010001", 23187 => "0110111110001010", 23188 => "0101010111000101", 23189 => "1110011000100010", 23190 => "0110011100011010", 23191 => "1010010001100110", 23192 => "0000111000010100", 23193 => "0100010110011111", 23194 => "1111111001100000", 23195 => "1000111110000010", 23196 => "1001111101011010", 23197 => "0010011010101011", 23198 => "0100110110010011", 23199 => "0010001111100111", 23200 => "1011101111101101", 23201 => "1001101011110010", 23202 => "1101100101110111", 23203 => "0011111110111001", 23204 => "0000101011111111", 23205 => "1110001100010001", 23206 => "0001000001101001", 23207 => "0000000111000111", 23208 => "1100000010001101", 23209 => "1001010100110110", 23210 => "1011001001001111", 23211 => "0010010010100101", 23212 => "1101001011000110", 23213 => "0000011101010111", 23214 => "0000100010001010", 23215 => "1010011100001111", 23216 => "1010101110011100", 23217 => "0011001001100011", 23218 => "0101010001110001", 23219 => "0111101101100001", 23220 => "0010101111001010", 23221 => "1000011101110101", 23222 => "0011100110010001", 23223 => "1100000110101111", 23224 => "1111111001000100", 23225 => "0000110111001110", 23226 => "1001011110010111", 23227 => "1111001100010011", 23228 => "1110110010100101", 23229 => "0110000011110001", 23230 => "1111010001110001", 23231 => "1110011010111001", 23232 => "0100001100101011", 23233 => "1100001100010101", 23234 => "0010001001000001", 23235 => "0000010110111000", 23236 => "0001001101001111", 23237 => "1000101010101110", 23238 => "0000001000001111", 23239 => "0001000110000001", 23240 => "1010101010010100", 23241 => "1100001101001001", 23242 => "0000111111000010", 23243 => "1100011010010010", 23244 => "0001100011111110", 23245 => "0111101111001111", 23246 => "1000010001010101", 23247 => "0010000101111010", 23248 => "1001000101110000", 23249 => "0011101001111111", 23250 => "0010000100000111", 23251 => "0101100001101101", 23252 => "1001000001010100", 23253 => "1001001111110001", 23254 => "1011100000010110", 23255 => "1111000110111111", 23256 => "0110111111000010", 23257 => "1101001100111010", 23258 => "0010100010110001", 23259 => "1010100011011001", 23260 => "0101101001101101", 23261 => "0011110110110110", 23262 => "1101110100000100", 23263 => "0001011011100110", 23264 => "1100110010000110", 23265 => "0110000101010101", 23266 => "1100101101000000", 23267 => "0100101000011010", 23268 => "0110000110011001", 23269 => "1111110000001110", 23270 => "0011001010011110", 23271 => "1101101100010100", 23272 => "0001110101101001", 23273 => "1101010001100010", 23274 => "1111100010100011", 23275 => "0111101111011011", 23276 => "1111011000110110", 23277 => "0111101101001110", 23278 => "0101010001101100", 23279 => "1110011010001111", 23280 => "1010011000111010", 23281 => "1000101110100100", 23282 => "1011011110100011", 23283 => "0010101010101100", 23284 => "1111101110001010", 23285 => "1010010100001111", 23286 => "0000000110100111", 23287 => "1101110010110010", 23288 => "0000100111001011", 23289 => "1001100011010100", 23290 => "1110010011011101", 23291 => "1111000110101001", 23292 => "1110111100111111", 23293 => "0110000100101001", 23294 => "0100101010101001", 23295 => "0010000111101010", 23296 => "0100001010011111", 23297 => "1100010111001010", 23298 => "0000011000001011", 23299 => "0101011010011100", 23300 => "0110101101011010", 23301 => "1110100011011110", 23302 => "1101001100101101", 23303 => "0100101001000111", 23304 => "0001011010011011", 23305 => "0010010101100101", 23306 => "0101001100101100", 23307 => "1101100100110011", 23308 => "0001110101010010", 23309 => "1000001111101101", 23310 => "1111100101011001", 23311 => "0101100000110010", 23312 => "1101101111010101", 23313 => "1001110100001101", 23314 => "0000101110110011", 23315 => "1011000000110000", 23316 => "1001000011100000", 23317 => "1011101001101011", 23318 => "0000111010001101", 23319 => "0001010000110011", 23320 => "1010010010010010", 23321 => "0001100010100001", 23322 => "1100111101111101", 23323 => "1101110011111010", 23324 => "1000010010000100", 23325 => "0001011000110100", 23326 => "0010111111100011", 23327 => "1100000101001000", 23328 => "0011000100100100", 23329 => "1111010100001011", 23330 => "0110010101101110", 23331 => "0011001101100110", 23332 => "0111111110111011", 23333 => "1000010001110111", 23334 => "1010011100100000", 23335 => "1100110001011000", 23336 => "1010100100011001", 23337 => "0010010110000001", 23338 => "1110101011110110", 23339 => "1111100101100010", 23340 => "1110101100000100", 23341 => "1110111101011110", 23342 => "1110001111110111", 23343 => "0111011110000000", 23344 => "1010111000000011", 23345 => "1001110010011000", 23346 => "0011110001010011", 23347 => "1111001100011101", 23348 => "0111001000101000", 23349 => "1111101000110001", 23350 => "0101110001101110", 23351 => "1101001101001001", 23352 => "1010000100100111", 23353 => "1100111011011110", 23354 => "1010001100111011", 23355 => "0110101101100010", 23356 => "1110111110110110", 23357 => "0100010011000011", 23358 => "1111100101110011", 23359 => "0011111101101011", 23360 => "0111010011011001", 23361 => "0011000000101110", 23362 => "0110111111101100", 23363 => "1000110110001000", 23364 => "1101100101001001", 23365 => "0100011000011010", 23366 => "0011100101000011", 23367 => "0000100010001010", 23368 => "1100001011010001", 23369 => "1011111000100011", 23370 => "0101110001101010", 23371 => "1110101111111100", 23372 => "1101000100100001", 23373 => "1111000110001000", 23374 => "0011101001000111", 23375 => "1110000100011001", 23376 => "1011111011011000", 23377 => "1111000011001101", 23378 => "0111011110110010", 23379 => "0101010101110100", 23380 => "0111100011011011", 23381 => "1011101011111010", 23382 => "0010100101111100", 23383 => "0111101101111010", 23384 => "0101101110000011", 23385 => "0000000100011001", 23386 => "1000100000011010", 23387 => "0110000100101010", 23388 => "1001011110111001", 23389 => "0010001100111000", 23390 => "0001000011101111", 23391 => "0110100010010001", 23392 => "0000100011111010", 23393 => "1111000000010110", 23394 => "1111101111110111", 23395 => "0000100001001110", 23396 => "0000110000100000", 23397 => "1010000001010010", 23398 => "1110011001010000", 23399 => "0100000010010101", 23400 => "1000000001101000", 23401 => "1000000101110010", 23402 => "1111001001001000", 23403 => "0000001110110100", 23404 => "1110011011011110", 23405 => "1111010001000001", 23406 => "0010001100010010", 23407 => "1011100010001101", 23408 => "1111111110011101", 23409 => "0001000011011101", 23410 => "1101101111100111", 23411 => "1101000011011010", 23412 => "1000111011001000", 23413 => "0000011111100010", 23414 => "1010110000111100", 23415 => "0111001101111100", 23416 => "1010100101100000", 23417 => "0100011010000001", 23418 => "1010111000011011", 23419 => "1010100010011011", 23420 => "1001011010110101", 23421 => "0010001011111100", 23422 => "1011010001111111", 23423 => "1001011000010100", 23424 => "0111101111101000", 23425 => "1001100010000111", 23426 => "1100010101001011", 23427 => "1001100110110110", 23428 => "1110011011110101", 23429 => "0000010010010011", 23430 => "1111110000011110", 23431 => "1010100010010101", 23432 => "1100111101011110", 23433 => "1100111111110110", 23434 => "1010011101101100", 23435 => "1001100000001000", 23436 => "1111011010000110", 23437 => "0101111000011110", 23438 => "1100100100101111", 23439 => "1001101011011001", 23440 => "1100110011110111", 23441 => "1010101111101011", 23442 => "0011010001001001", 23443 => "0001101111101011", 23444 => "0000010111101111", 23445 => "1101000101000000", 23446 => "0000011011010010", 23447 => "1110001111010110", 23448 => "0011100000010000", 23449 => "1101101010001001", 23450 => "0001010111100010", 23451 => "0000010100100000", 23452 => "0101101101000001", 23453 => "1100010111101000", 23454 => "0001101000011110", 23455 => "0111000010101010", 23456 => "0011010000111110", 23457 => "0110001011010111", 23458 => "1011010100111000", 23459 => "0011100011110011", 23460 => "0111111010111010", 23461 => "1011101110001111", 23462 => "0001101100001100", 23463 => "0101011110011101", 23464 => "0111010111000111", 23465 => "1011100100111000", 23466 => "1010000111011110", 23467 => "1001111101101111", 23468 => "0110100001101101", 23469 => "1001011110111001", 23470 => "0010000110010001", 23471 => "1010000010110111", 23472 => "0000110100111011", 23473 => "1111101110010111", 23474 => "1011110010101100", 23475 => "0000100110010010", 23476 => "0100101000011001", 23477 => "0000001001001101", 23478 => "1010001110010000", 23479 => "1001001000010011", 23480 => "0000000010101001", 23481 => "0001110000111100", 23482 => "0000011100011111", 23483 => "0111011111001101", 23484 => "1010010011101111", 23485 => "0000001010100010", 23486 => "0001101111111001", 23487 => "1100011100001100", 23488 => "1011111111000100", 23489 => "0101010110101011", 23490 => "0110010100001101", 23491 => "0111011000101010", 23492 => "1110001101110000", 23493 => "0100010110011110", 23494 => "1001010100110010", 23495 => "0000001011010011", 23496 => "0111101101100011", 23497 => "1000000000101111", 23498 => "1110011011101101", 23499 => "0101100101100101", 23500 => "0100110110101111", 23501 => "1101100010001100", 23502 => "1110110010001011", 23503 => "0011101111010010", 23504 => "0111110000111011", 23505 => "1100111110000101", 23506 => "0101110110001010", 23507 => "1100000011110101", 23508 => "0001000000101010", 23509 => "0111000010111110", 23510 => "1010100101100101", 23511 => "1011011110101110", 23512 => "1010100100001001", 23513 => "0100011110101110", 23514 => "0010110101101010", 23515 => "1100011101000010", 23516 => "1111110010100101", 23517 => "1001001101101010", 23518 => "0001010100011111", 23519 => "0000010111111001", 23520 => "0111001011001010", 23521 => "0101001011000100", 23522 => "0111111100010000", 23523 => "1100100100001010", 23524 => "0100011011000110", 23525 => "1011110110011011", 23526 => "1110000000110100", 23527 => "0011100000000000", 23528 => "0010111010001010", 23529 => "0100011110011100", 23530 => "0000011011110110", 23531 => "0011001000011100", 23532 => "1011011110011000", 23533 => "1110011100101111", 23534 => "1100101110111100", 23535 => "0000001111100110", 23536 => "1000100110001011", 23537 => "0101010100100001", 23538 => "0011110101000101", 23539 => "0000010100000000", 23540 => "1111110110001001", 23541 => "1110110101111010", 23542 => "1100100000000101", 23543 => "1000111111101001", 23544 => "1011001000010011", 23545 => "0011001111100000", 23546 => "1111110101000110", 23547 => "0110110011110110", 23548 => "0110111101111001", 23549 => "1100011100001110", 23550 => "1110010000111010", 23551 => "0001010001010110", 23552 => "1110001100000101", 23553 => "1011000010101110", 23554 => "0110001101010010", 23555 => "0001100111100110", 23556 => "1111000101100101", 23557 => "0000000000001101", 23558 => "0100010001011010", 23559 => "0101100001001001", 23560 => "1011001100010011", 23561 => "1000011101110001", 23562 => "0000010100000000", 23563 => "0101000101101111", 23564 => "1111101110000001", 23565 => "0111010111110011", 23566 => "0010100111101111", 23567 => "1010111010010100", 23568 => "0011110000011011", 23569 => "0001010111111111", 23570 => "0101101000110111", 23571 => "0010011001100010", 23572 => "0011010000010110", 23573 => "0100001000100111", 23574 => "0000010101111011", 23575 => "0001100010001111", 23576 => "0100101010111111", 23577 => "1100001000101110", 23578 => "1110000101101111", 23579 => "0011001100010000", 23580 => "1101010101110110", 23581 => "0110011100100110", 23582 => "0101010110010100", 23583 => "0010001111110100", 23584 => "0010011101100001", 23585 => "0001110111101011", 23586 => "0000100010011100", 23587 => "1011110111011110", 23588 => "1100001010101111", 23589 => "0111001110011110", 23590 => "1110111101100001", 23591 => "0111011101111011", 23592 => "0001110101001100", 23593 => "1001000001000100", 23594 => "0011000010011001", 23595 => "0101100111011011", 23596 => "1110111000111000", 23597 => "1010100011000011", 23598 => "0111101110001010", 23599 => "1010100010110100", 23600 => "0000010100101000", 23601 => "1010011100001110", 23602 => "0110110100111000", 23603 => "0011001000010111", 23604 => "0001101001101011", 23605 => "1101010111001000", 23606 => "0001100110011100", 23607 => "0000110100011111", 23608 => "1101001101111111", 23609 => "0000010000010010", 23610 => "0010111101000101", 23611 => "1000001100110101", 23612 => "0001011001001100", 23613 => "0100100010001010", 23614 => "0010001001001110", 23615 => "0101010111010001", 23616 => "0000001001010100", 23617 => "1111111000101100", 23618 => "0110011110001101", 23619 => "1110111111111010", 23620 => "0100000010111100", 23621 => "0011011110010101", 23622 => "0001001011110010", 23623 => "1010011001010100", 23624 => "0000100110000000", 23625 => "1100100010111010", 23626 => "1101010101110100", 23627 => "0010010111101110", 23628 => "0001000001101011", 23629 => "1011110001001000", 23630 => "1001000011001110", 23631 => "1101101111001101", 23632 => "1010110010010100", 23633 => "0100000110010011", 23634 => "1111010011100010", 23635 => "0000111000011101", 23636 => "1110001110000111", 23637 => "1010111001111000", 23638 => "0011100100011000", 23639 => "1011000001010010", 23640 => "1011100110100101", 23641 => "0010001011111110", 23642 => "0101000101100011", 23643 => "1011001001101101", 23644 => "0101111001110001", 23645 => "0010010010000001", 23646 => "0011110100000101", 23647 => "0011010001101101", 23648 => "1101111111101011", 23649 => "0001011000101101", 23650 => "0111101100000101", 23651 => "1110101000101101", 23652 => "1111110101101110", 23653 => "1101111010110001", 23654 => "1001100001101111", 23655 => "1100110011111011", 23656 => "0001110111101111", 23657 => "0100101001111110", 23658 => "1101011001000100", 23659 => "1001101110110110", 23660 => "1010101001101101", 23661 => "1000001001111010", 23662 => "0010001011110010", 23663 => "0011001100010111", 23664 => "0101111111100100", 23665 => "0101000011000000", 23666 => "1111010000100011", 23667 => "0010010111100010", 23668 => "1001011001101001", 23669 => "0010100000100010", 23670 => "0110110100001111", 23671 => "1000001110111100", 23672 => "1000111111010000", 23673 => "0100000101100011", 23674 => "1010001011001110", 23675 => "0111111101011010", 23676 => "1001100101111010", 23677 => "0111011100110101", 23678 => "1110000001001000", 23679 => "0010010000110011", 23680 => "0000110000010000", 23681 => "1000110101110110", 23682 => "0010110100000101", 23683 => "0010111011010000", 23684 => "1110001110011110", 23685 => "0001111101110100", 23686 => "1100000001111110", 23687 => "0001000110000110", 23688 => "1001001011100101", 23689 => "0001001100110100", 23690 => "1110000000000010", 23691 => "0100010000011000", 23692 => "1111001101110011", 23693 => "1011001011011010", 23694 => "0111000000101110", 23695 => "1011010100001001", 23696 => "1000100110100100", 23697 => "1100010111010100", 23698 => "0001100000110001", 23699 => "0001000011011110", 23700 => "0000111111111111", 23701 => "0011100001001010", 23702 => "1110111100010001", 23703 => "0110011001000011", 23704 => "1110010010111010", 23705 => "0101100000110111", 23706 => "0010000011101010", 23707 => "1011100011000101", 23708 => "0001110111100011", 23709 => "0011111011001011", 23710 => "1111010100011001", 23711 => "0101101011111111", 23712 => "1011010100001110", 23713 => "1100110111101110", 23714 => "0100011110011101", 23715 => "0100111000001101", 23716 => "0111000011101110", 23717 => "1101001100110001", 23718 => "0011000100100101", 23719 => "0000111011010111", 23720 => "1110101110110111", 23721 => "0011101010010110", 23722 => "0011011101010110", 23723 => "0011110010010011", 23724 => "0001111010110111", 23725 => "1000010001000101", 23726 => "0000011101001000", 23727 => "1000111001100010", 23728 => "0011101111001100", 23729 => "0000000110001100", 23730 => "0110010110010000", 23731 => "1110111001001010", 23732 => "0010010110000011", 23733 => "0011000100100000", 23734 => "1010000100111000", 23735 => "0111011101001110", 23736 => "0011100100001000", 23737 => "0010010101010011", 23738 => "1101001101101100", 23739 => "1010111100100111", 23740 => "0100000100110101", 23741 => "0010011001111110", 23742 => "1101100011011100", 23743 => "0101101100100001", 23744 => "0101000011111110", 23745 => "0000011111010001", 23746 => "1110111101100010", 23747 => "0110101001101011", 23748 => "1100111011111010", 23749 => "0011010011000111", 23750 => "0110011101111110", 23751 => "1001000001000101", 23752 => "1010101000100010", 23753 => "1001110110110100", 23754 => "1110001111010011", 23755 => "1100010100110110", 23756 => "1010111111011101", 23757 => "1001000110011010", 23758 => "0011101111101110", 23759 => "1111100101000010", 23760 => "1011101110110110", 23761 => "1011101101110000", 23762 => "0011000101111001", 23763 => "0011010100100111", 23764 => "1100001111000100", 23765 => "1011000100010101", 23766 => "0010110011100000", 23767 => "0011101011001000", 23768 => "0010001101110001", 23769 => "0011001000101001", 23770 => "0100011010100111", 23771 => "0101100011111010", 23772 => "0100110111001101", 23773 => "1110001000100110", 23774 => "0111000110100100", 23775 => "0110101110111101", 23776 => "1100010100001110", 23777 => "0011001000100010", 23778 => "1001011010110100", 23779 => "1110000100110011", 23780 => "1111001011011100", 23781 => "0000110011010011", 23782 => "1001001010101100", 23783 => "1010110001110001", 23784 => "1110001011100011", 23785 => "0000100101011001", 23786 => "1011110000000010", 23787 => "0011110100001101", 23788 => "0001011111000011", 23789 => "1110000100111101", 23790 => "0011001010001101", 23791 => "1000001100110101", 23792 => "1101011100100101", 23793 => "1010110100101101", 23794 => "0000110101110111", 23795 => "0001110000111110", 23796 => "0010010101011111", 23797 => "1100001111010100", 23798 => "1101110011101010", 23799 => "1101001110111110", 23800 => "0101010100110111", 23801 => "0001110001101000", 23802 => "0101010001000001", 23803 => "0101000111000111", 23804 => "0001110101111001", 23805 => "0010111010110111", 23806 => "1010010101000101", 23807 => "0011010110011100", 23808 => "0101001111010011", 23809 => "1000001011011111", 23810 => "0000110000110011", 23811 => "0000001011110000", 23812 => "1101000111101010", 23813 => "0011100100101010", 23814 => "1100101001001001", 23815 => "1010110100100001", 23816 => "0110100011111010", 23817 => "1001110100100010", 23818 => "0001001111011101", 23819 => "0001010100110011", 23820 => "1110000101000110", 23821 => "0010001011011010", 23822 => "0110111110100111", 23823 => "1110111010110010", 23824 => "1111110101101011", 23825 => "1011111011101111", 23826 => "1111100110111001", 23827 => "0100000000000111", 23828 => "1000110111011110", 23829 => "1000011011001001", 23830 => "0111010100001110", 23831 => "1111110110010010", 23832 => "0111110111110100", 23833 => "0101000100011010", 23834 => "0111100010101001", 23835 => "0111000001011000", 23836 => "1000001101101001", 23837 => "1101101001101001", 23838 => "0000011101010100", 23839 => "1010001110001101", 23840 => "0000111100011011", 23841 => "0000101010010000", 23842 => "1000011010110001", 23843 => "1110001110000100", 23844 => "0011100010101100", 23845 => "0001000101001101", 23846 => "0101011001000101", 23847 => "1011100100111100", 23848 => "0100101010111011", 23849 => "0100101000001100", 23850 => "0000111101100100", 23851 => "0010100011111010", 23852 => "0001010101110101", 23853 => "0100100100011011", 23854 => "0011010000011000", 23855 => "1000010011111000", 23856 => "1111101011000101", 23857 => "0100010001011111", 23858 => "1100111101101010", 23859 => "1010100101001010", 23860 => "0110000101000101", 23861 => "0100010100011101", 23862 => "0001111110011010", 23863 => "0010100110100110", 23864 => "1101110000001100", 23865 => "1110000100100010", 23866 => "1100111100010110", 23867 => "1100111110100100", 23868 => "1000000001010010", 23869 => "0000001011010000", 23870 => "1010100100111010", 23871 => "1100010111110011", 23872 => "0111111101000001", 23873 => "1100110010111110", 23874 => "0110001001001011", 23875 => "0011111000100000", 23876 => "1111000101001000", 23877 => "1001111011111010", 23878 => "0100101100011000", 23879 => "0001011111000100", 23880 => "0100111000001011", 23881 => "1111000100111111", 23882 => "0000101001100110", 23883 => "0110001101101111", 23884 => "1001110011000110", 23885 => "0011011101001010", 23886 => "1000011010000110", 23887 => "1100100010100100", 23888 => "0000001111011011", 23889 => "0101010011001111", 23890 => "0111010001101011", 23891 => "0111011011010111", 23892 => "0101111001101101", 23893 => "1010111110010101", 23894 => "1111111100110111", 23895 => "1101101100000101", 23896 => "0011000100111100", 23897 => "0101101100000010", 23898 => "0101111001000001", 23899 => "0111101000001011", 23900 => "0101011111110001", 23901 => "1110011111110101", 23902 => "1000101010111100", 23903 => "0110001110111101", 23904 => "0111111000110100", 23905 => "1001001110001101", 23906 => "1010111101101110", 23907 => "0011110000100111", 23908 => "0100101100100111", 23909 => "1110111101010010", 23910 => "1010001111111011", 23911 => "1110111110111100", 23912 => "0111001001001111", 23913 => "1100011110110010", 23914 => "0101100100011010", 23915 => "0011000011001000", 23916 => "0110010001101111", 23917 => "0000110010001111", 23918 => "1011101011001000", 23919 => "1010100100010101", 23920 => "1110101011001000", 23921 => "1000011101001000", 23922 => "0110010000010111", 23923 => "1011110100011111", 23924 => "0001000010110001", 23925 => "0101101110101011", 23926 => "0000101101000111", 23927 => "1100110101110100", 23928 => "0010000010010011", 23929 => "0110100011110101", 23930 => "1010000101011100", 23931 => "0101011000110000", 23932 => "1001010010010101", 23933 => "1110010110100110", 23934 => "0011010100011010", 23935 => "0100110111100100", 23936 => "1101000011000011", 23937 => "1100000000101000", 23938 => "1010001001110000", 23939 => "0001011010100000", 23940 => "1111111100101110", 23941 => "0010101011100111", 23942 => "1011100000100100", 23943 => "1001110111110101", 23944 => "0100011100111000", 23945 => "0101110111011011", 23946 => "0101100011010000", 23947 => "1010100011010001", 23948 => "0001010011001000", 23949 => "0101110001100001", 23950 => "0001011001011100", 23951 => "1010000011111110", 23952 => "0110111001100111", 23953 => "1100011101000001", 23954 => "1110010101111011", 23955 => "1011000011010000", 23956 => "0110010101010010", 23957 => "1111100100101000", 23958 => "1111010111100010", 23959 => "1110110110101101", 23960 => "0111101101110000", 23961 => "1111101001010011", 23962 => "0111010000111111", 23963 => "1111111000101110", 23964 => "1111010100101100", 23965 => "1101100111110111", 23966 => "1111011111100101", 23967 => "0110111100101001", 23968 => "1110110011110100", 23969 => "1101000010101010", 23970 => "1010011001111100", 23971 => "1101010100001000", 23972 => "0000011001111101", 23973 => "0110010100110110", 23974 => "1011001000101111", 23975 => "0100011111001111", 23976 => "0111000101100011", 23977 => "0011111010000110", 23978 => "0101001011001101", 23979 => "0011100000011011", 23980 => "1001100000111111", 23981 => "0111100011001110", 23982 => "0011100110101010", 23983 => "1011011101111111", 23984 => "1010101010010011", 23985 => "1011110000110101", 23986 => "0001000000000010", 23987 => "1010010111110111", 23988 => "0011001000100110", 23989 => "1100000111000010", 23990 => "0010011100111101", 23991 => "1000100011000001", 23992 => "0011010010101011", 23993 => "1110111001111011", 23994 => "0100000101011101", 23995 => "0000111101011101", 23996 => "1110010110010010", 23997 => "1010101010111000", 23998 => "0111110100000001", 23999 => "1111010001100111", 24000 => "0101001011101001", 24001 => "0010110000101101", 24002 => "0011001001010101", 24003 => "1001111111101100", 24004 => "1010011100011000", 24005 => "1111111011001011", 24006 => "0101101000100011", 24007 => "1110110101000000", 24008 => "1000001101111000", 24009 => "1000000010101000", 24010 => "1110111101001000", 24011 => "0011101101101000", 24012 => "1111001111010100", 24013 => "0000000111010001", 24014 => "1000111011001111", 24015 => "0101010110001000", 24016 => "0111011011100001", 24017 => "0100110011010110", 24018 => "0101000101010110", 24019 => "1010000101100110", 24020 => "1000111010001101", 24021 => "1011010001001100", 24022 => "1011110101000011", 24023 => "0110101100000011", 24024 => "0101010001101100", 24025 => "0110100100000101", 24026 => "0011000101011010", 24027 => "1010100111101011", 24028 => "0110000101101100", 24029 => "0001001001001011", 24030 => "1001101001100100", 24031 => "0011101110010111", 24032 => "0001111101101000", 24033 => "0111000101110000", 24034 => "0110010010110001", 24035 => "0001011010100101", 24036 => "0101111001111001", 24037 => "0010000101011100", 24038 => "0111100101100101", 24039 => "1100100000001000", 24040 => "1001100101101101", 24041 => "0010001011111101", 24042 => "0011110010101101", 24043 => "0011111110110111", 24044 => "1010010100110000", 24045 => "0100000100110010", 24046 => "0101100110001100", 24047 => "1010001010000000", 24048 => "1100100110101010", 24049 => "0111111011011011", 24050 => "1111100111111000", 24051 => "0110000001111101", 24052 => "0011000101011001", 24053 => "1100111001000101", 24054 => "0000110100100001", 24055 => "1111010100111000", 24056 => "0110110000110010", 24057 => "0110101011100010", 24058 => "1101011100011101", 24059 => "0001100010110111", 24060 => "1011111011000100", 24061 => "0001111100101001", 24062 => "1011100100110101", 24063 => "1000100100111100", 24064 => "0110010100001101", 24065 => "0110001100101101", 24066 => "0110001010001000", 24067 => "0000000001011000", 24068 => "1110100100110000", 24069 => "0000011100001100", 24070 => "0100011111100110", 24071 => "0111110111110011", 24072 => "0001110000011010", 24073 => "0110000100100111", 24074 => "1101101011010111", 24075 => "1010100101100011", 24076 => "1011001000011010", 24077 => "1100101110111010", 24078 => "0111100010001001", 24079 => "0011000001010110", 24080 => "0011001100011010", 24081 => "1110101000011010", 24082 => "1111110000110011", 24083 => "0000100100010001", 24084 => "0001100001010111", 24085 => "0011010000100011", 24086 => "1011110101001000", 24087 => "1110111101101011", 24088 => "0110011000010001", 24089 => "1000110000100100", 24090 => "0000001110101001", 24091 => "1011100001100011", 24092 => "0000010110001010", 24093 => "1111101110101100", 24094 => "0111000111010011", 24095 => "0111100010101110", 24096 => "0010010100101001", 24097 => "0100100100110011", 24098 => "0000001011001111", 24099 => "0101001001010110", 24100 => "1000110101101000", 24101 => "1001000111000001", 24102 => "0110111011111011", 24103 => "0001100111110000", 24104 => "0011101110110110", 24105 => "1101000001111111", 24106 => "1100111011010011", 24107 => "0011010101010001", 24108 => "1011101100110011", 24109 => "0100101000110010", 24110 => "0010111000101100", 24111 => "1010110100101111", 24112 => "0111000110111101", 24113 => "1101010101100000", 24114 => "1110101100010100", 24115 => "0011110000001111", 24116 => "1101101101000110", 24117 => "0010101101011111", 24118 => "1111001011110111", 24119 => "1110100100100110", 24120 => "1010000010111000", 24121 => "0010111110100010", 24122 => "1111001000100110", 24123 => "1000111110100011", 24124 => "0000110001001110", 24125 => "1101110000111101", 24126 => "1010000011110101", 24127 => "0010100110000110", 24128 => "1111110111111011", 24129 => "0010001000010110", 24130 => "0011000110100100", 24131 => "0011000101001111", 24132 => "1010000000111001", 24133 => "0000001111100100", 24134 => "0110110000100111", 24135 => "1110100001101011", 24136 => "0101001001100011", 24137 => "1010011111111100", 24138 => "0110000000100100", 24139 => "0101010110111011", 24140 => "1111111000101011", 24141 => "0111110100111101", 24142 => "0110100101011110", 24143 => "0000000000101110", 24144 => "0110011000010001", 24145 => "0011000000111011", 24146 => "1100110111010010", 24147 => "1000111010111101", 24148 => "1000111110100111", 24149 => "0010000001111110", 24150 => "1111101110000011", 24151 => "0101011101000001", 24152 => "0100000101101010", 24153 => "1001101101110101", 24154 => "1010100110001101", 24155 => "1000010001101101", 24156 => "0100110001101111", 24157 => "1000110001010101", 24158 => "1111001000010111", 24159 => "0110011011001011", 24160 => "1011010100001110", 24161 => "1111011110001101", 24162 => "0010101100100101", 24163 => "1100111001100000", 24164 => "1011011000011010", 24165 => "0000010011011000", 24166 => "0101001100100110", 24167 => "0101000010011001", 24168 => "1010010010001101", 24169 => "0100001011100110", 24170 => "0000000100011000", 24171 => "0100110010010011", 24172 => "1101001101110101", 24173 => "0111101001001100", 24174 => "0000110101101010", 24175 => "0101110100101101", 24176 => "0011000011110111", 24177 => "1001111110100101", 24178 => "1000110010011000", 24179 => "1010000100111100", 24180 => "1110110100001001", 24181 => "0001000001110001", 24182 => "1100111111110010", 24183 => "1001010100000011", 24184 => "0101011101111001", 24185 => "1101111110101101", 24186 => "0001000101001000", 24187 => "1110111011101000", 24188 => "0111111010101111", 24189 => "0011010010100111", 24190 => "1010100001011011", 24191 => "0001110011111111", 24192 => "0011000111110100", 24193 => "1111001110110011", 24194 => "1011111001100000", 24195 => "0100110110001010", 24196 => "1010101110011010", 24197 => "1011101001101000", 24198 => "1011100110000111", 24199 => "0001010101111010", 24200 => "1010011101010101", 24201 => "0111011011001010", 24202 => "1011000100011010", 24203 => "1111110011011101", 24204 => "1001110011100101", 24205 => "0001001110101101", 24206 => "0001000011111110", 24207 => "1011010111000100", 24208 => "0111001101010010", 24209 => "1011100001010101", 24210 => "1001101010101101", 24211 => "0100101011111110", 24212 => "1010110111011111", 24213 => "1100101111110101", 24214 => "1000100110110001", 24215 => "0100000011101101", 24216 => "1011100011010111", 24217 => "0011111010101111", 24218 => "1101101010000000", 24219 => "0111111100000110", 24220 => "1001000100010101", 24221 => "1111100100111101", 24222 => "1110000001111000", 24223 => "1011000001101011", 24224 => "1101001101101001", 24225 => "0011100000111000", 24226 => "1100101101000011", 24227 => "0110101001000101", 24228 => "1000001011001011", 24229 => "1010011100101100", 24230 => "0111010111001010", 24231 => "0111111101001000", 24232 => "1101011001100001", 24233 => "0011100001110101", 24234 => "1001000011011001", 24235 => "0101111010110101", 24236 => "1111000101101011", 24237 => "1111110100010011", 24238 => "1001100010011011", 24239 => "0000111100101010", 24240 => "0010010101010000", 24241 => "0101000111000110", 24242 => "1000100000011001", 24243 => "0000010010111011", 24244 => "1011000000110101", 24245 => "0011101010111001", 24246 => "0000010000110000", 24247 => "1001000001100000", 24248 => "0000101011111011", 24249 => "1001110111001011", 24250 => "0000111000011001", 24251 => "1100010101001011", 24252 => "1000110101101010", 24253 => "0101100111001001", 24254 => "0001110011101001", 24255 => "1010001101000100", 24256 => "1101000000111110", 24257 => "1101111101110011", 24258 => "1000110010010000", 24259 => "1010111010001011", 24260 => "0000010100110100", 24261 => "0101011001111110", 24262 => "1001111011111000", 24263 => "1001110101110001", 24264 => "0111010011100011", 24265 => "1011011010101001", 24266 => "0100011100110000", 24267 => "1011100000000011", 24268 => "1010100011101100", 24269 => "1100100101001111", 24270 => "1010101000100101", 24271 => "1011100010010010", 24272 => "0110011011001011", 24273 => "1110001111111000", 24274 => "0011010000100101", 24275 => "1110000010100000", 24276 => "0001100001000100", 24277 => "0110111110010011", 24278 => "1100101010111100", 24279 => "0011110101011101", 24280 => "0100101101101001", 24281 => "0111111100111000", 24282 => "0101111101110100", 24283 => "0101001101010100", 24284 => "1011001011110111", 24285 => "1001101100000111", 24286 => "0101011000110100", 24287 => "1011011100110011", 24288 => "1000000000111100", 24289 => "0011010100000110", 24290 => "1000010101101110", 24291 => "1010100111100101", 24292 => "0011101110110001", 24293 => "0001101010110111", 24294 => "0111111111101000", 24295 => "1001111001000111", 24296 => "0100110011110101", 24297 => "1011101000011001", 24298 => "0100011101001011", 24299 => "1001010101011000", 24300 => "0000000101110111", 24301 => "1010101000001101", 24302 => "1111100001110101", 24303 => "0111011110000110", 24304 => "1011111011001101", 24305 => "0000001111110100", 24306 => "0100010000110011", 24307 => "1111010010101011", 24308 => "0111101001111010", 24309 => "0011000010110010", 24310 => "1000100100001111", 24311 => "1011110001001001", 24312 => "1010101101101100", 24313 => "0101110100010000", 24314 => "1100100110001110", 24315 => "1000100000001001", 24316 => "0110011100001100", 24317 => "1000111111100100", 24318 => "1110000010010011", 24319 => "0001001110101000", 24320 => "0010111011010000", 24321 => "1101101010111110", 24322 => "0101001000010110", 24323 => "0010100100111001", 24324 => "1100000111000011", 24325 => "1001010111100100", 24326 => "0011001001110100", 24327 => "1111100000010000", 24328 => "1100110001110111", 24329 => "1111111101010010", 24330 => "1011000110000101", 24331 => "1000101000011001", 24332 => "1011100011110111", 24333 => "1101010001010110", 24334 => "1101100100010000", 24335 => "0110010110000110", 24336 => "0101001101000101", 24337 => "0101011001101010", 24338 => "0011010001100100", 24339 => "1110111111111110", 24340 => "1001111100001100", 24341 => "0110111000100100", 24342 => "0011101000001000", 24343 => "1110001010110110", 24344 => "1010000110010000", 24345 => "0101111101110010", 24346 => "0000011100111001", 24347 => "0011111100100101", 24348 => "1100100111100011", 24349 => "0001111010100110", 24350 => "1011011110011110", 24351 => "1100000011111100", 24352 => "0100100000101111", 24353 => "0000001101000001", 24354 => "0110100100001010", 24355 => "1100000011101011", 24356 => "1010111011111101", 24357 => "0101110010011001", 24358 => "1111000101100110", 24359 => "1001001000010011", 24360 => "0100011110010100", 24361 => "1100010100010100", 24362 => "0101000110111001", 24363 => "1111111101110000", 24364 => "1011000100010111", 24365 => "1101100011001000", 24366 => "1001111010010011", 24367 => "1011001111010000", 24368 => "0010111101010011", 24369 => "0100100000110010", 24370 => "0010001110110101", 24371 => "0001010101101101", 24372 => "0001000111110101", 24373 => "1110110010110111", 24374 => "0110000001010000", 24375 => "1101111111111111", 24376 => "0110110100010111", 24377 => "1011111100011010", 24378 => "1111000010010101", 24379 => "0001111011100010", 24380 => "0011001001001001", 24381 => "0111110111101100", 24382 => "0001001011010010", 24383 => "1011001100110000", 24384 => "1011100101111011", 24385 => "0001010110110011", 24386 => "0111100010111000", 24387 => "0100100101011110", 24388 => "1100110011101101", 24389 => "1110111101010011", 24390 => "1110010001110001", 24391 => "0100011111010100", 24392 => "0110101110011100", 24393 => "0111001110100000", 24394 => "0010100100001111", 24395 => "1111101100101101", 24396 => "1000111001000111", 24397 => "1001001100111110", 24398 => "1100100101100010", 24399 => "0100110110101011", 24400 => "1110010000101100", 24401 => "0101100101000101", 24402 => "1101110001010011", 24403 => "1011000101110111", 24404 => "0101001111111001", 24405 => "1011100000010001", 24406 => "1001001000111000", 24407 => "1101011000110010", 24408 => "1011001000011100", 24409 => "0110011010110011", 24410 => "0110001101110100", 24411 => "1010001010110010", 24412 => "1101101111010111", 24413 => "1110101100000000", 24414 => "1110010011001110", 24415 => "1101010011101010", 24416 => "0111111101110110", 24417 => "0001000001000011", 24418 => "0011111011000010", 24419 => "0100111110001101", 24420 => "1011110011110100", 24421 => "0110000101011111", 24422 => "0111111001101000", 24423 => "1111100001100011", 24424 => "0110010000111100", 24425 => "0011001000110010", 24426 => "0011110011000110", 24427 => "0101101100010000", 24428 => "0000010100100110", 24429 => "1011101010011100", 24430 => "0001001010010011", 24431 => "1101000110110001", 24432 => "0101110100000001", 24433 => "0011011001110100", 24434 => "0110111101110010", 24435 => "0111011101101100", 24436 => "0101100101001100", 24437 => "0000001100100011", 24438 => "1111101110111110", 24439 => "1100000000000011", 24440 => "0101010011011110", 24441 => "1010011011001010", 24442 => "0000000111101100", 24443 => "1010111011110111", 24444 => "0100001001011000", 24445 => "0101000011101110", 24446 => "1001101101101111", 24447 => "1010001001110100", 24448 => "1001000000101011", 24449 => "1011010101001110", 24450 => "0101011011010101", 24451 => "0000010010111011", 24452 => "0011010111000010", 24453 => "0010001001111100", 24454 => "1000011011001000", 24455 => "1111101110000111", 24456 => "0100001100101111", 24457 => "0100000010110011", 24458 => "0100111100010001", 24459 => "0101001100011111", 24460 => "0011110010101110", 24461 => "0011001100111011", 24462 => "1101001011101111", 24463 => "1101011110100000", 24464 => "0110110011010011", 24465 => "0100101001010001", 24466 => "0100111000000101", 24467 => "0111001110010111", 24468 => "0110010111001100", 24469 => "1101001011101011", 24470 => "1000101111011100", 24471 => "0110000101111111", 24472 => "0000100101110100", 24473 => "1001000010001000", 24474 => "0100000000010010", 24475 => "0111010100011111", 24476 => "0111010010111100", 24477 => "0111001000010100", 24478 => "0101000101111000", 24479 => "0001010100110101", 24480 => "1110001010010000", 24481 => "1101100010100111", 24482 => "0010110111101111", 24483 => "1111111101110010", 24484 => "0101000011101011", 24485 => "0000110110001100", 24486 => "1000110100000000", 24487 => "0001111110010101", 24488 => "1000011001001110", 24489 => "0111101001111110", 24490 => "1001010101010110", 24491 => "0001100101011000", 24492 => "1011010100111101", 24493 => "0110110100110111", 24494 => "1101111110011111", 24495 => "0000111010001001", 24496 => "0111110011110111", 24497 => "1110100111101111", 24498 => "0000011010110101", 24499 => "1001000000101111", 24500 => "0010001111001011", 24501 => "1111101100111000", 24502 => "0000010101010101", 24503 => "1101111001101001", 24504 => "1100100011011010", 24505 => "0011000101001001", 24506 => "0010110111101111", 24507 => "1001010111011101", 24508 => "1010001110111111", 24509 => "0100101100101000", 24510 => "1101101000010100", 24511 => "0100011011010010", 24512 => "0111111100000111", 24513 => "0001101110011101", 24514 => "1000011001011000", 24515 => "0000110110010000", 24516 => "0101010101011111", 24517 => "0000100001100000", 24518 => "1101010101000000", 24519 => "0001011010001110", 24520 => "0001110111110001", 24521 => "0000001101011100", 24522 => "1100111010001111", 24523 => "0000111011011100", 24524 => "1111101010011110", 24525 => "1000001011111100", 24526 => "1010111010110010", 24527 => "0011110101110000", 24528 => "0111000011100001", 24529 => "1101010001111101", 24530 => "1111111100001101", 24531 => "1100101000111110", 24532 => "1010011001001010", 24533 => "0110101111010010", 24534 => "0011011101010010", 24535 => "1101110010100100", 24536 => "0111111101001010", 24537 => "0010110001011110", 24538 => "0001111110111010", 24539 => "0010111101010010", 24540 => "0011111000010010", 24541 => "1110110110100000", 24542 => "1010010010000010", 24543 => "1101110101000110", 24544 => "1110101100010011", 24545 => "0100010011001000", 24546 => "0110111100101011", 24547 => "1100101111110100", 24548 => "1001101111110100", 24549 => "0011111001011000", 24550 => "1001001111111100", 24551 => "1110010101100101", 24552 => "0011001111001000", 24553 => "1111111111010000", 24554 => "0001101011101010", 24555 => "0000010111111101", 24556 => "1110100000011001", 24557 => "0001101111111000", 24558 => "1100111110000111", 24559 => "0000110001011001", 24560 => "1110010101101110", 24561 => "1100111011110100", 24562 => "1001010100101110", 24563 => "1000101000100011", 24564 => "1110010010001100", 24565 => "1000011001011110", 24566 => "0101010111001000", 24567 => "1011000010001101", 24568 => "0101010111100101", 24569 => "0111001011010000", 24570 => "0111000010101111", 24571 => "1111111000000000", 24572 => "1001011011101110", 24573 => "0110100000000000", 24574 => "1010000111000010", 24575 => "1110011101011011", 24576 => "1001110100001001", 24577 => "0000110001101011", 24578 => "1110000011100100", 24579 => "0001111010100010", 24580 => "1101111000100000", 24581 => "1111100010110111", 24582 => "1110100111110011", 24583 => "1101101100001111", 24584 => "0100110111100101", 24585 => "0010111011010101", 24586 => "0110101101000000", 24587 => "0001010001010111", 24588 => "1010001101111110", 24589 => "0110110011000101", 24590 => "0001000101111101", 24591 => "0100011101000001", 24592 => "0100010100011111", 24593 => "0101011000001100", 24594 => "0110000101100101", 24595 => "1101000110001100", 24596 => "1010111010000011", 24597 => "0000100001101111", 24598 => "0101100001001000", 24599 => "0100010101101110", 24600 => "0100001011000001", 24601 => "1001000000001111", 24602 => "0101010011011000", 24603 => "1111110111001010", 24604 => "0111111001100000", 24605 => "1111100010101110", 24606 => "1000000000000000", 24607 => "0111101101100001", 24608 => "1001000111001001", 24609 => "1010000011010100", 24610 => "1001111010111000", 24611 => "0001000000001000", 24612 => "0111100010101110", 24613 => "0010000001101100", 24614 => "1101110000101110", 24615 => "0110000000111001", 24616 => "1010010110100010", 24617 => "0110110010100100", 24618 => "1111011111010111", 24619 => "0001111000111010", 24620 => "0111111110000101", 24621 => "1001000010011111", 24622 => "1110110110011111", 24623 => "0011101101001111", 24624 => "0010100111001100", 24625 => "1011100101110011", 24626 => "1000110011000011", 24627 => "1110101111011111", 24628 => "1100100010011000", 24629 => "0101000111100110", 24630 => "1000111001010000", 24631 => "1101001001101101", 24632 => "0110001010001100", 24633 => "0101001011011000", 24634 => "1100000011000000", 24635 => "0100000101011100", 24636 => "1010111100010110", 24637 => "1101000000001001", 24638 => "1000001100101100", 24639 => "1111111010101110", 24640 => "1001001001111010", 24641 => "0111111100110011", 24642 => "0110011110011001", 24643 => "0001100001111011", 24644 => "0100011101110111", 24645 => "1000001001100100", 24646 => "0110000110111111", 24647 => "1110110011110001", 24648 => "0011111111101000", 24649 => "0010101010100110", 24650 => "0100110000010011", 24651 => "1011011000011011", 24652 => "1011001011001110", 24653 => "0011101100111010", 24654 => "0011011110101100", 24655 => "0110110111100000", 24656 => "1101010100000100", 24657 => "0010101011101011", 24658 => "0101000111100101", 24659 => "1011000110011110", 24660 => "0001000100100111", 24661 => "0000001000001111", 24662 => "0000010111011001", 24663 => "1101011011010101", 24664 => "1101010011100100", 24665 => "0110001010011001", 24666 => "0110001000110110", 24667 => "0011010010110111", 24668 => "1100101001111010", 24669 => "1101100011000111", 24670 => "1001111011111000", 24671 => "1011000111100110", 24672 => "0001100110110111", 24673 => "1101100101001000", 24674 => "1110110111100100", 24675 => "1011111000111010", 24676 => "1011001110100010", 24677 => "1000001100111010", 24678 => "0110000000011110", 24679 => "1000110010100100", 24680 => "0001111111110001", 24681 => "1101110010101111", 24682 => "1011010101011011", 24683 => "1110111101110000", 24684 => "0001100101001001", 24685 => "1000001001111001", 24686 => "0111001001001001", 24687 => "1001011100101111", 24688 => "0101000110100011", 24689 => "0001101000100110", 24690 => "1000001011010010", 24691 => "0110110001000001", 24692 => "0011101001011011", 24693 => "1110011001011100", 24694 => "1100111111110111", 24695 => "0001111010001111", 24696 => "0100110101110101", 24697 => "0101000010001011", 24698 => "1011110101101111", 24699 => "0111100011110111", 24700 => "0000010001110110", 24701 => "1001100010000010", 24702 => "0111111001111101", 24703 => "0100111100000010", 24704 => "1110001111110111", 24705 => "0101101001111001", 24706 => "0100110000100110", 24707 => "0101000010110110", 24708 => "0111101100001101", 24709 => "1000101100101100", 24710 => "1001111111100111", 24711 => "1001110010110000", 24712 => "1011010100100110", 24713 => "0001111001010100", 24714 => "0000011001010001", 24715 => "1010100111010000", 24716 => "1100011011101010", 24717 => "0001101001111010", 24718 => "0100111100011111", 24719 => "1110011010001010", 24720 => "1001011110100000", 24721 => "0101000101000101", 24722 => "0011101101101110", 24723 => "0001001101000001", 24724 => "1011000101110101", 24725 => "0111000010001110", 24726 => "1010001110001110", 24727 => "0111010101111010", 24728 => "0011110001111000", 24729 => "1000110111110111", 24730 => "0010010100100110", 24731 => "1011001000110101", 24732 => "0101111000001110", 24733 => "1000000100010110", 24734 => "0001100111110010", 24735 => "1010110011111101", 24736 => "1001011101010001", 24737 => "1000010100111101", 24738 => "1100000000111010", 24739 => "0110101100111011", 24740 => "1010001001110011", 24741 => "0111100111110101", 24742 => "1101100010010100", 24743 => "1001000011001100", 24744 => "0101110001010101", 24745 => "1000101010101000", 24746 => "0010110010111011", 24747 => "0111000111110101", 24748 => "0110011001010010", 24749 => "1010010011100000", 24750 => "1001101001010001", 24751 => "0100011101010001", 24752 => "0010000000110000", 24753 => "0110110100011101", 24754 => "0111100011110000", 24755 => "0100001011011101", 24756 => "0010101101000101", 24757 => "0011000101101100", 24758 => "1100111010110101", 24759 => "1110110110010111", 24760 => "1111011111111111", 24761 => "1100110100000011", 24762 => "0011110111010010", 24763 => "1101011110011110", 24764 => "1011100101001000", 24765 => "0100011111001001", 24766 => "0111010001010110", 24767 => "0000000011100100", 24768 => "0110100101111100", 24769 => "1011101001100000", 24770 => "0111101101001101", 24771 => "1001000101011000", 24772 => "1001010010110010", 24773 => "1111100011000001", 24774 => "0000001001001000", 24775 => "1111010011010110", 24776 => "1010000010110110", 24777 => "0100000110010011", 24778 => "1101000010111000", 24779 => "1010010101110000", 24780 => "1111111110100001", 24781 => "0110001011000100", 24782 => "1110101100100011", 24783 => "0010100000101111", 24784 => "0111101010110000", 24785 => "1101111110101100", 24786 => "0110010010000000", 24787 => "1110100011101100", 24788 => "0100101011001100", 24789 => "0111101100001110", 24790 => "1111011111111011", 24791 => "1011001101000000", 24792 => "1111011100110101", 24793 => "0110011110000011", 24794 => "0101101111001010", 24795 => "0000111011011000", 24796 => "1010000101110000", 24797 => "0010110101101010", 24798 => "1111000110011110", 24799 => "1101111011111100", 24800 => "1010010100001100", 24801 => "0010011111010110", 24802 => "1100100011111110", 24803 => "0110011111011100", 24804 => "0111000101100110", 24805 => "1010100010000011", 24806 => "1111011111110101", 24807 => "1000101011000100", 24808 => "0100100001000111", 24809 => "0011001010001100", 24810 => "1001110101011110", 24811 => "0000110011001010", 24812 => "1100100110110000", 24813 => "0000000100000001", 24814 => "1100000001000101", 24815 => "0110111101101010", 24816 => "0000110010011001", 24817 => "0001000110110011", 24818 => "0101100100100010", 24819 => "0000100001100010", 24820 => "0000100110000101", 24821 => "0100000100001010", 24822 => "0111001010001010", 24823 => "1000011111100110", 24824 => "0111111010001001", 24825 => "1001011001001000", 24826 => "0110110110001000", 24827 => "0011011011011110", 24828 => "0101110001110011", 24829 => "1111001100011110", 24830 => "1111100011100110", 24831 => "1101110111010000", 24832 => "1101111111011101", 24833 => "1100100000100000", 24834 => "0101000010111000", 24835 => "1111100001011001", 24836 => "1001000011000000", 24837 => "0010010101001100", 24838 => "1101111110010010", 24839 => "1111100100010001", 24840 => "1010110111011101", 24841 => "1001010010001100", 24842 => "0001101110010101", 24843 => "1011101011010010", 24844 => "1100001001100111", 24845 => "1111101111100001", 24846 => "1001000110011000", 24847 => "0101001000100011", 24848 => "0111111011100001", 24849 => "0110011001001101", 24850 => "1110110000100110", 24851 => "1111100110000011", 24852 => "1111101000101010", 24853 => "0011110001000111", 24854 => "0000001010000110", 24855 => "1001011000001100", 24856 => "0100100101110101", 24857 => "1010010001111110", 24858 => "0110100111111111", 24859 => "0001100100111110", 24860 => "1111101110110000", 24861 => "0101100011110011", 24862 => "1000001010010000", 24863 => "1111101110011100", 24864 => "0011010111110110", 24865 => "0101001010111000", 24866 => "1011011100011111", 24867 => "1011101010010101", 24868 => "0100000001111000", 24869 => "0001011010110101", 24870 => "0100111001101111", 24871 => "1010101011110001", 24872 => "1011000100001110", 24873 => "1011110011110010", 24874 => "1111010110011010", 24875 => "0000011000001101", 24876 => "0100011001100000", 24877 => "0011010110000110", 24878 => "1111001101000110", 24879 => "1111111011100011", 24880 => "1110011001001000", 24881 => "0110100000111111", 24882 => "0111011101010101", 24883 => "1100100001011110", 24884 => "0100011001110110", 24885 => "0001111010010111", 24886 => "0101100100001110", 24887 => "1101010010111001", 24888 => "1100011001011010", 24889 => "0000101001101101", 24890 => "1111010001110110", 24891 => "1001011011101011", 24892 => "1010010001010001", 24893 => "1111110111101000", 24894 => "1101001100111000", 24895 => "0110100001101110", 24896 => "0101110011111101", 24897 => "1010111111100111", 24898 => "0011001110010110", 24899 => "0111100001011001", 24900 => "1011100110000001", 24901 => "1001110011001011", 24902 => "1110100011001111", 24903 => "1010000000110110", 24904 => "1111100100000000", 24905 => "1110110010111011", 24906 => "1010001010100010", 24907 => "1010011111011100", 24908 => "1101011010000110", 24909 => "1110010011101100", 24910 => "1010101010000111", 24911 => "0011000010010000", 24912 => "0010101101000100", 24913 => "1101100110010111", 24914 => "1001101110001011", 24915 => "1101110110101110", 24916 => "0100110001011100", 24917 => "1010010110100100", 24918 => "1000111100100011", 24919 => "1000100101101000", 24920 => "0100111100111100", 24921 => "0000010100010101", 24922 => "0111011111101001", 24923 => "0111001001100110", 24924 => "0110010111011010", 24925 => "1111010110100011", 24926 => "0110100101101110", 24927 => "0100000111011001", 24928 => "1011001110101101", 24929 => "0110000001001110", 24930 => "0001100010011001", 24931 => "0111011100101101", 24932 => "0100110101001100", 24933 => "1011100011110001", 24934 => "0111110010000111", 24935 => "0001011110110001", 24936 => "1010100110100010", 24937 => "0011000011111100", 24938 => "1010101101001000", 24939 => "1101111000011010", 24940 => "1001100111001111", 24941 => "1000111111001000", 24942 => "1000110111001100", 24943 => "0010011001001100", 24944 => "0000100100111010", 24945 => "1111011000010110", 24946 => "1001001010011011", 24947 => "1101001011010000", 24948 => "1001001001010101", 24949 => "0010101100000011", 24950 => "0110001110011111", 24951 => "1101110001111011", 24952 => "0110011000111011", 24953 => "0101010110010010", 24954 => "1100111011001010", 24955 => "1011010010011010", 24956 => "1001000010010011", 24957 => "0110101010111111", 24958 => "1011011100001011", 24959 => "1101100001110101", 24960 => "0101000110111101", 24961 => "0110000001001001", 24962 => "0010001110110011", 24963 => "1110000110000100", 24964 => "1110010010111100", 24965 => "0000110011000010", 24966 => "1011010111011011", 24967 => "0011101010110000", 24968 => "0000010010000101", 24969 => "1001100110010011", 24970 => "0011111010111100", 24971 => "1100110011110010", 24972 => "1101111110001100", 24973 => "1001110000011011", 24974 => "0001011011100101", 24975 => "0010101100011110", 24976 => "1000111011011011", 24977 => "0110011110011101", 24978 => "0101100101010010", 24979 => "1100001111001110", 24980 => "1001010100101101", 24981 => "1101111100110110", 24982 => "0000110001010011", 24983 => "1110101101011101", 24984 => "0101111010101010", 24985 => "0011010000010111", 24986 => "1101100111101010", 24987 => "1101000010000001", 24988 => "0111100001111000", 24989 => "1011001001110111", 24990 => "0111100000011001", 24991 => "1101000001101010", 24992 => "0011011011010111", 24993 => "1110110111101101", 24994 => "1000101000110010", 24995 => "1111101001000101", 24996 => "1000010100101010", 24997 => "0011001000101011", 24998 => "1011010000001100", 24999 => "1001101011000010", 25000 => "1111001111000010", 25001 => "1111110010100101", 25002 => "1100111110100001", 25003 => "1110010011001000", 25004 => "0001010111110011", 25005 => "0000101010000110", 25006 => "0110100000001001", 25007 => "0111000110000100", 25008 => "0010111101011101", 25009 => "1011001110111000", 25010 => "0000110000110001", 25011 => "1111111010100001", 25012 => "1101110100100111", 25013 => "1111110000111101", 25014 => "0000010001011000", 25015 => "1101111110101101", 25016 => "1001000011110101", 25017 => "1110110010000000", 25018 => "1010001010000001", 25019 => "1011101001000000", 25020 => "0001111100011110", 25021 => "0101100110111001", 25022 => "1110000011101001", 25023 => "0101001101010100", 25024 => "0011001001011101", 25025 => "1100110011101010", 25026 => "1100111101101010", 25027 => "0001111101101110", 25028 => "0010111101101100", 25029 => "1100011010101111", 25030 => "1110100110101001", 25031 => "0000010101010101", 25032 => "0101010110001110", 25033 => "0110101101000001", 25034 => "0110111011011000", 25035 => "0101111000010111", 25036 => "1010111110111000", 25037 => "1001001010111110", 25038 => "1010100010001101", 25039 => "1111100100010010", 25040 => "1001001110110010", 25041 => "1000000011000111", 25042 => "0011111101101111", 25043 => "0110111100100010", 25044 => "1100011110011011", 25045 => "0101001110010111", 25046 => "1111110010111110", 25047 => "1110000111001110", 25048 => "1100101011011001", 25049 => "1001011100101000", 25050 => "1101110000110011", 25051 => "1110100001000001", 25052 => "1100101001010010", 25053 => "1110100011001010", 25054 => "1001011100010001", 25055 => "1111101101000000", 25056 => "1100110000011011", 25057 => "1110010100111001", 25058 => "1101111010010110", 25059 => "1110001011010011", 25060 => "0000100011000111", 25061 => "1111100000011001", 25062 => "1110010001101101", 25063 => "1000101011111111", 25064 => "1110000011001001", 25065 => "0010111111110101", 25066 => "0010001111010000", 25067 => "1000011100111000", 25068 => "1110000111011000", 25069 => "1010100111101111", 25070 => "1101100110010110", 25071 => "0000010000111001", 25072 => "1001101100010111", 25073 => "0000011000000111", 25074 => "1111110011110001", 25075 => "1110110010011010", 25076 => "1101111011010101", 25077 => "0110010101110101", 25078 => "1010010011011111", 25079 => "1111010001000011", 25080 => "0100110010000010", 25081 => "0100100101100100", 25082 => "0100110101110110", 25083 => "0011100011011111", 25084 => "0101110001100100", 25085 => "1001101111110010", 25086 => "1111010000001011", 25087 => "0011101011000100", 25088 => "0001010000000100", 25089 => "1111110000101011", 25090 => "1011000100000001", 25091 => "1111000100010000", 25092 => "1101110111010001", 25093 => "1000010101110010", 25094 => "1101111100101111", 25095 => "1101100100010110", 25096 => "0111111001001001", 25097 => "1001110011101010", 25098 => "0000111010111000", 25099 => "1001010001001100", 25100 => "0000110101000100", 25101 => "1101011100111010", 25102 => "0111111001101101", 25103 => "1000100101100000", 25104 => "1100000001111011", 25105 => "0111100111110100", 25106 => "1101011111101111", 25107 => "0111011011011000", 25108 => "0001011010010110", 25109 => "0000011100001101", 25110 => "0000111010011110", 25111 => "1001010100111001", 25112 => "1000010011011110", 25113 => "1011011111011001", 25114 => "1100100000001101", 25115 => "0110111101100010", 25116 => "1000101110110100", 25117 => "1111001001101001", 25118 => "1111101101001101", 25119 => "1000011110101111", 25120 => "1110001000001100", 25121 => "0011001001011000", 25122 => "1101110110001000", 25123 => "0111110110111011", 25124 => "1001011000011010", 25125 => "1110110101001101", 25126 => "0001011100110000", 25127 => "0101110101110000", 25128 => "0000011011101010", 25129 => "0010111100101010", 25130 => "1110011101001001", 25131 => "1101111011100011", 25132 => "0101111010000011", 25133 => "0100000010001010", 25134 => "1010111010110001", 25135 => "1000010110010011", 25136 => "0111100011110101", 25137 => "1000010110000111", 25138 => "0111011010010001", 25139 => "1101000000101101", 25140 => "1110001000000001", 25141 => "1010111110001001", 25142 => "0001000000000000", 25143 => "1010010011011001", 25144 => "1100011101111101", 25145 => "0010011111100101", 25146 => "0000010101111010", 25147 => "1010110100101110", 25148 => "1110100110110101", 25149 => "1001100101011101", 25150 => "1000100110110011", 25151 => "1111010110000111", 25152 => "1001011101001011", 25153 => "0011010100101110", 25154 => "0010010011001010", 25155 => "1100100011110011", 25156 => "0101010011000001", 25157 => "0011100101100100", 25158 => "0111100011110111", 25159 => "0111011100001111", 25160 => "1010100111100101", 25161 => "1011000111101110", 25162 => "0111110100101111", 25163 => "0101101010001110", 25164 => "0100100001011010", 25165 => "0001101101100110", 25166 => "0000011111001000", 25167 => "1100001000110010", 25168 => "0101001011100011", 25169 => "1111011010110000", 25170 => "0100000110000100", 25171 => "0011010001111111", 25172 => "0111101011001110", 25173 => "0101100010110100", 25174 => "0000001000110010", 25175 => "0010111100001001", 25176 => "1001110100010100", 25177 => "0101111000111100", 25178 => "0100110000010010", 25179 => "0100011000110101", 25180 => "0011110011001100", 25181 => "0001000010111000", 25182 => "0101110011111010", 25183 => "1000010100101100", 25184 => "0011100000011111", 25185 => "0001111110100011", 25186 => "1100011011000100", 25187 => "0000001100101110", 25188 => "1001110110010000", 25189 => "1011011111011100", 25190 => "0100101101100001", 25191 => "0000101011111011", 25192 => "0110111110100110", 25193 => "1111001111010101", 25194 => "1100000000010101", 25195 => "0100011010000101", 25196 => "0001111011001011", 25197 => "1100100101101100", 25198 => "0001111000101001", 25199 => "0101111111110010", 25200 => "1011011100010101", 25201 => "0110100000110011", 25202 => "1000100010111111", 25203 => "0010001001001100", 25204 => "1000010000101011", 25205 => "0111101011011100", 25206 => "0010111110011011", 25207 => "0100110111010111", 25208 => "0011011101111111", 25209 => "0101001110011000", 25210 => "1000001001110101", 25211 => "0111100000001100", 25212 => "0111101000111100", 25213 => "1000001110101011", 25214 => "0101100010101100", 25215 => "1011001111100000", 25216 => "1110001101001111", 25217 => "0111100110011111", 25218 => "1100000011110111", 25219 => "1010011101110101", 25220 => "0011000111011011", 25221 => "0000010011001101", 25222 => "0111100001100001", 25223 => "1010110100001000", 25224 => "0010010110011111", 25225 => "0011010101111000", 25226 => "1100100011111011", 25227 => "1001100000111110", 25228 => "1100011001010011", 25229 => "0110100110110101", 25230 => "0110011010100100", 25231 => "1111011100010001", 25232 => "0011101001000101", 25233 => "1001000001011101", 25234 => "1101100010010110", 25235 => "1011100001011100", 25236 => "1010001000010110", 25237 => "0101001000010110", 25238 => "1010000110010111", 25239 => "0001011001011001", 25240 => "1000101000010001", 25241 => "0101010000010101", 25242 => "1101011010101010", 25243 => "0101110110111001", 25244 => "0101110000001111", 25245 => "0101010001010011", 25246 => "1011111000011101", 25247 => "1101101010000000", 25248 => "1100111100011000", 25249 => "0001011111001100", 25250 => "1001101011010110", 25251 => "0110010000010101", 25252 => "0011111011011110", 25253 => "0000101111110100", 25254 => "1110110001101110", 25255 => "0101001010100111", 25256 => "1011100110011100", 25257 => "0001010110010101", 25258 => "0101110101110001", 25259 => "0111100110100011", 25260 => "1110010110001100", 25261 => "0011011100000111", 25262 => "1011010010101101", 25263 => "0000110110001010", 25264 => "1101001001101111", 25265 => "1100100011100100", 25266 => "0110111111010100", 25267 => "0100011011001010", 25268 => "0101000101011110", 25269 => "1010111001010111", 25270 => "0101100101001000", 25271 => "1001110001100000", 25272 => "0000000001101110", 25273 => "1001001001101111", 25274 => "0101110111000011", 25275 => "0011010001011010", 25276 => "1111110100100001", 25277 => "0001001100101100", 25278 => "0101110000100100", 25279 => "1100001100111000", 25280 => "0111001001110111", 25281 => "1100000001011100", 25282 => "0001011011000011", 25283 => "1011011000011001", 25284 => "0101001100110011", 25285 => "1101010110011101", 25286 => "0011000111010101", 25287 => "1110000100011011", 25288 => "1101110001000001", 25289 => "0111001001010011", 25290 => "1011101110110111", 25291 => "1110111011100110", 25292 => "1001101110101001", 25293 => "1100111000100101", 25294 => "0110000100011101", 25295 => "0110000110010100", 25296 => "0000011000010100", 25297 => "0010000010101011", 25298 => "1010111101100100", 25299 => "0010001011110101", 25300 => "1001001110001101", 25301 => "1000000011110100", 25302 => "0000100110010100", 25303 => "0111010011011011", 25304 => "1110101001011010", 25305 => "0100001101010110", 25306 => "1011001100110001", 25307 => "1011100100010100", 25308 => "1001001011011011", 25309 => "1011111111011010", 25310 => "1010010101000000", 25311 => "1101001011000111", 25312 => "0101110011010011", 25313 => "1100000101000111", 25314 => "1100110111011001", 25315 => "1111101111011010", 25316 => "0010010001100110", 25317 => "1001101101000001", 25318 => "1000001111111000", 25319 => "0000111011010001", 25320 => "0001100011100110", 25321 => "1101111100101001", 25322 => "1001100000001100", 25323 => "0111001011010000", 25324 => "1001001001111011", 25325 => "1001111101101010", 25326 => "1010100100100101", 25327 => "1001010001000010", 25328 => "0111010010110111", 25329 => "0110110111101010", 25330 => "1011100011100111", 25331 => "1010110010000110", 25332 => "0010101011011111", 25333 => "0101110111000001", 25334 => "0111000101110100", 25335 => "1111100101010011", 25336 => "1100101010011110", 25337 => "1010110110001011", 25338 => "1110000110000111", 25339 => "1011001100110001", 25340 => "0110011101110010", 25341 => "1001010110111101", 25342 => "0110110001001111", 25343 => "0001110110101011", 25344 => "0000111101101001", 25345 => "0000111010110010", 25346 => "1011101000110100", 25347 => "0110110111010000", 25348 => "1001110101101111", 25349 => "1001011010001010", 25350 => "0110111001100011", 25351 => "0110011111100111", 25352 => "1011111000111101", 25353 => "1000100101000101", 25354 => "1101001011101000", 25355 => "1010001011001100", 25356 => "1010110011001100", 25357 => "1011011000101010", 25358 => "1010110011110010", 25359 => "1101101101001111", 25360 => "1011101011010111", 25361 => "0011100101010111", 25362 => "0011100011110011", 25363 => "0111111010001011", 25364 => "1101011010100100", 25365 => "1100100010000010", 25366 => "0110100111100010", 25367 => "0001000000101000", 25368 => "0100110001010100", 25369 => "0000000001100101", 25370 => "1010111110101000", 25371 => "1010000011000111", 25372 => "1010110111000000", 25373 => "1011110100100011", 25374 => "0001000011001111", 25375 => "1110001001111100", 25376 => "0111000011011011", 25377 => "0110010100010010", 25378 => "0011110100101001", 25379 => "0001000111011011", 25380 => "0011000001001110", 25381 => "1011111111001110", 25382 => "0100001111000110", 25383 => "0001111011000010", 25384 => "1100010010000111", 25385 => "0001011110111100", 25386 => "0011001000111000", 25387 => "0011010001100100", 25388 => "0010001100000000", 25389 => "0011111000110100", 25390 => "1111111010010100", 25391 => "0010100110101101", 25392 => "0110111110011101", 25393 => "0101100100010000", 25394 => "0110100100100111", 25395 => "0001010110001010", 25396 => "1111111000110100", 25397 => "1010110010100011", 25398 => "1011101111100001", 25399 => "0111000000010101", 25400 => "0101101001110101", 25401 => "1110111011101011", 25402 => "1100000000010011", 25403 => "0011110001000010", 25404 => "1000011010100100", 25405 => "1111010000011101", 25406 => "1111001001100111", 25407 => "1100110111100001", 25408 => "0010000001011001", 25409 => "0011100011010111", 25410 => "0100111011100100", 25411 => "0110111101111001", 25412 => "0100001110111011", 25413 => "0111100101001110", 25414 => "0001101011110000", 25415 => "0011001110101001", 25416 => "1001110000010011", 25417 => "0110111000111110", 25418 => "1010001001001000", 25419 => "1101110101010111", 25420 => "0010001100101011", 25421 => "0000001101101101", 25422 => "0110111011101001", 25423 => "0111010010111001", 25424 => "1000010111011010", 25425 => "0001101001110100", 25426 => "1011111001001100", 25427 => "1100010111111110", 25428 => "1101011101010011", 25429 => "1100100001110011", 25430 => "0000111010101101", 25431 => "0111110001011111", 25432 => "1111000110000100", 25433 => "1110000001110110", 25434 => "1110101000010111", 25435 => "1100001001011111", 25436 => "1110100010110001", 25437 => "1000011010010010", 25438 => "0111100010001011", 25439 => "1101011011111111", 25440 => "0000010001101011", 25441 => "0010010101101010", 25442 => "1110100111001100", 25443 => "0010010010101110", 25444 => "0100111111101000", 25445 => "1011011011001101", 25446 => "0010011011010101", 25447 => "1110110110110111", 25448 => "1111011011110101", 25449 => "1111010101011111", 25450 => "0111110100110100", 25451 => "1001111010100001", 25452 => "1000110100011101", 25453 => "1110011010101111", 25454 => "0010011110011100", 25455 => "1110011000111010", 25456 => "0011000101010100", 25457 => "0101010000001011", 25458 => "0110110101000110", 25459 => "1000110111100101", 25460 => "1001110101101000", 25461 => "0110111111101110", 25462 => "1110010101111111", 25463 => "1001010101110001", 25464 => "1001001000010010", 25465 => "0001100100101110", 25466 => "1111010100011111", 25467 => "1011110011000000", 25468 => "0111110010110110", 25469 => "0100010111111101", 25470 => "1101010011001001", 25471 => "0011000001011110", 25472 => "0010110010000101", 25473 => "1000110011101110", 25474 => "1011101010000101", 25475 => "0001101101110110", 25476 => "1011111001011100", 25477 => "1111110010111111", 25478 => "1011111111100000", 25479 => "1010000101111100", 25480 => "0100110100110000", 25481 => "0100100101010110", 25482 => "0100000011000110", 25483 => "0001010100111101", 25484 => "1011111110111000", 25485 => "0011101101100000", 25486 => "1010110000010011", 25487 => "0001101101000101", 25488 => "1010110001110010", 25489 => "0101101010011100", 25490 => "0101101111000000", 25491 => "0001000001000100", 25492 => "0010110100100011", 25493 => "1000011011001010", 25494 => "0010101001011000", 25495 => "1000110110111101", 25496 => "1111010000100000", 25497 => "1001011100011101", 25498 => "0111001100011110", 25499 => "1001100011000101", 25500 => "1110101100110100", 25501 => "1110000010100111", 25502 => "1101011101110001", 25503 => "1101011000101111", 25504 => "0000100111110111", 25505 => "1010101100011101", 25506 => "1100000000010011", 25507 => "1001000101000010", 25508 => "0001000110100010", 25509 => "1000101010111111", 25510 => "0110111011101001", 25511 => "1001010111100101", 25512 => "0010101010010101", 25513 => "0100001010111011", 25514 => "1011111111001000", 25515 => "1110011011100111", 25516 => "1101110011101010", 25517 => "0110011000100010", 25518 => "1010111000101101", 25519 => "1011101111011110", 25520 => "1011001011001101", 25521 => "1010000110101111", 25522 => "1100011110000110", 25523 => "0000000001111000", 25524 => "1111110000100101", 25525 => "1111010101101010", 25526 => "0000001000110110", 25527 => "1100001101001100", 25528 => "1101000011111101", 25529 => "0001011101011111", 25530 => "0101000011000010", 25531 => "0101000110100110", 25532 => "1111000101100010", 25533 => "0110100111111111", 25534 => "1010101100000011", 25535 => "1001101011110100", 25536 => "1101000010000111", 25537 => "1101000001011011", 25538 => "0111100110011011", 25539 => "1001101111001011", 25540 => "0011001100010111", 25541 => "0011010111010100", 25542 => "0010000010000101", 25543 => "0100101011100010", 25544 => "0010000110101110", 25545 => "0000001111100110", 25546 => "1100010001101100", 25547 => "1110101001111010", 25548 => "1110101111101011", 25549 => "1100000110000101", 25550 => "0000010111100100", 25551 => "1010000100001100", 25552 => "0111110001100011", 25553 => "1100010010010011", 25554 => "0001000110000000", 25555 => "1110101111010001", 25556 => "0110111001000010", 25557 => "0111100010111010", 25558 => "1100101010110010", 25559 => "0100100101110010", 25560 => "0011100101010001", 25561 => "0001000111000011", 25562 => "1011100000010100", 25563 => "1110101110111001", 25564 => "1110000011000010", 25565 => "0010000010110010", 25566 => "0111000000111100", 25567 => "1001000101001101", 25568 => "0111011101110011", 25569 => "1100101001100101", 25570 => "1011101111100011", 25571 => "1100001111011100", 25572 => "0101110111011110", 25573 => "1101001101011010", 25574 => "0000011101101011", 25575 => "1111010001000001", 25576 => "1100011011001110", 25577 => "0010110100011100", 25578 => "1001100101111110", 25579 => "0011101110110111", 25580 => "1010011101110111", 25581 => "0011111100110011", 25582 => "1101001001111000", 25583 => "0110110101110001", 25584 => "1000101010010010", 25585 => "0101011111011010", 25586 => "1010011111100000", 25587 => "1010110110110110", 25588 => "0010110110110011", 25589 => "1001011101001001", 25590 => "0100101000100000", 25591 => "1110001011010111", 25592 => "1011000011011101", 25593 => "1001111001110110", 25594 => "1011001010101111", 25595 => "1011111010100000", 25596 => "1010001111010010", 25597 => "0101000111000111", 25598 => "0011001111101111", 25599 => "1100011111011001", 25600 => "0110111000111010", 25601 => "0111001000010100", 25602 => "1010000111011101", 25603 => "0001010010001001", 25604 => "0100000000110100", 25605 => "0111100110100110", 25606 => "0110111000011100", 25607 => "0100110010001110", 25608 => "1010010001010111", 25609 => "0101111011011101", 25610 => "1100001010100001", 25611 => "0111011100000101", 25612 => "1100101000001010", 25613 => "1010101100000001", 25614 => "0001011110110111", 25615 => "0101011010011000", 25616 => "1111100100101010", 25617 => "1101001100101101", 25618 => "0000010100000000", 25619 => "0000101101110111", 25620 => "1010100111100101", 25621 => "0101110101111000", 25622 => "1101100111010101", 25623 => "1000100100001010", 25624 => "1101010100100111", 25625 => "1010010100101110", 25626 => "0011000011011110", 25627 => "0101011100100101", 25628 => "0111011001001011", 25629 => "1011000011010010", 25630 => "0011011111010100", 25631 => "1101111100110011", 25632 => "1101011111001001", 25633 => "0101101111011000", 25634 => "1011101000110001", 25635 => "1011001011001011", 25636 => "0110111100001010", 25637 => "0001111000111010", 25638 => "1100001101100010", 25639 => "0101001001011000", 25640 => "1101001110100011", 25641 => "0010111010010000", 25642 => "1101001110010010", 25643 => "1110000100111101", 25644 => "1000001111100101", 25645 => "0000000000100001", 25646 => "0101111000111000", 25647 => "1011110110110101", 25648 => "1111100101111111", 25649 => "0100110001101101", 25650 => "0100100101110101", 25651 => "1101011010110000", 25652 => "0110101110100010", 25653 => "0001001111101011", 25654 => "1101001110001111", 25655 => "1000001100101110", 25656 => "0101001110011101", 25657 => "1010101011011110", 25658 => "1100111110111001", 25659 => "0001010100010110", 25660 => "0010011011000000", 25661 => "1111100101100000", 25662 => "0010011010011110", 25663 => "0100110101001001", 25664 => "0110001000100111", 25665 => "0101011001100110", 25666 => "0101011100000000", 25667 => "0110001000011110", 25668 => "1001111011100001", 25669 => "1111011100110010", 25670 => "1011000010100101", 25671 => "0000010100001001", 25672 => "1001110000100110", 25673 => "0110101100010111", 25674 => "0100010111101101", 25675 => "0010101011011110", 25676 => "0100010101011101", 25677 => "1000001110010101", 25678 => "1111110010010101", 25679 => "0001001011000111", 25680 => "1101111001001100", 25681 => "1011110010001011", 25682 => "0101001000101100", 25683 => "0101010001100010", 25684 => "1000001011011100", 25685 => "1101111100000110", 25686 => "1001011010100111", 25687 => "0100101101011011", 25688 => "1011101011011110", 25689 => "0010001001001111", 25690 => "0110110001000011", 25691 => "1100110010011010", 25692 => "1101011001000100", 25693 => "1110110101000010", 25694 => "0010001100100110", 25695 => "0001100110010010", 25696 => "0110111011001011", 25697 => "1110001111010110", 25698 => "1000011010000000", 25699 => "1010100100110000", 25700 => "0100001010111100", 25701 => "0010111010110001", 25702 => "0011110010000110", 25703 => "1100011001010100", 25704 => "1110100000111011", 25705 => "0010110110110011", 25706 => "0000110101111110", 25707 => "0001101000011011", 25708 => "0110000010000011", 25709 => "1110101011110000", 25710 => "1101111011010011", 25711 => "1110000000000000", 25712 => "1110111001111111", 25713 => "1100010100011001", 25714 => "0110110100111100", 25715 => "1111100010011000", 25716 => "0101110111001110", 25717 => "1001100000100011", 25718 => "1000101010010000", 25719 => "0110000000001000", 25720 => "1111100001100011", 25721 => "1111100100111101", 25722 => "0011101001001110", 25723 => "1111010111000111", 25724 => "1110010010011011", 25725 => "0011010000001011", 25726 => "0001010010100110", 25727 => "1000101101111001", 25728 => "0111001101100101", 25729 => "1000100101001001", 25730 => "0010111010001101", 25731 => "0101110101100101", 25732 => "1100010101001111", 25733 => "0010010100111110", 25734 => "0111101000011100", 25735 => "0101010011010001", 25736 => "0001011101001110", 25737 => "1010101101001110", 25738 => "1100001101100000", 25739 => "0111101000001110", 25740 => "0001110001001101", 25741 => "1010110111101101", 25742 => "0111111101011001", 25743 => "0001101010101000", 25744 => "1111000010000111", 25745 => "1010100000111111", 25746 => "0101011001111110", 25747 => "0111001011100100", 25748 => "1000001111110000", 25749 => "0111101101000010", 25750 => "0100100110001100", 25751 => "0011000110011001", 25752 => "1101010100100110", 25753 => "0011011010111111", 25754 => "1110001010110100", 25755 => "0011011111111111", 25756 => "1010101101100100", 25757 => "0000011101000101", 25758 => "0011000100000101", 25759 => "1000100101010111", 25760 => "1011000110100010", 25761 => "0110010110010110", 25762 => "0011111001001110", 25763 => "1001010010100100", 25764 => "0011011101000001", 25765 => "0100000000000101", 25766 => "0001011101000010", 25767 => "1000011110000100", 25768 => "1010101000011111", 25769 => "0110110110010101", 25770 => "1111101010111101", 25771 => "0010011101011100", 25772 => "0111000110010010", 25773 => "0110110010001101", 25774 => "1111111110000101", 25775 => "1000110000010011", 25776 => "0101001110100110", 25777 => "0101010000101111", 25778 => "0000001001010111", 25779 => "1010111111000110", 25780 => "1000010110011010", 25781 => "0000000011101000", 25782 => "1100011010101001", 25783 => "0100110000011010", 25784 => "1111111111100110", 25785 => "1001000110011001", 25786 => "1001011100000110", 25787 => "0001101011000000", 25788 => "0011010000110100", 25789 => "1110101101000111", 25790 => "0010011000111010", 25791 => "0101011100000000", 25792 => "1001011010100111", 25793 => "0110100111111010", 25794 => "1101010101110010", 25795 => "0001000000101100", 25796 => "1100111110000011", 25797 => "0000101101111111", 25798 => "0100111110001100", 25799 => "0010111010010011", 25800 => "1010001011010001", 25801 => "0100101111010011", 25802 => "0100000011111010", 25803 => "0100000111101000", 25804 => "1100011001000011", 25805 => "1000110011100001", 25806 => "0000101110101111", 25807 => "1110001110101100", 25808 => "0011011001111000", 25809 => "0000110010110001", 25810 => "1100001011100011", 25811 => "1001100100011111", 25812 => "0001101111111011", 25813 => "1110101100110100", 25814 => "1101001101011111", 25815 => "0111010100011001", 25816 => "0010000101101010", 25817 => "1111101111101100", 25818 => "1001111111100000", 25819 => "1001101000010101", 25820 => "1010101101100111", 25821 => "0010001001001001", 25822 => "1011010011011000", 25823 => "1100001001110100", 25824 => "0100011000110010", 25825 => "0010111001100101", 25826 => "0100000001001110", 25827 => "1100001101010011", 25828 => "1001011011010000", 25829 => "1110011100101011", 25830 => "0011100001111010", 25831 => "1101001100100001", 25832 => "0110000000001011", 25833 => "1110011101111110", 25834 => "0110000110110001", 25835 => "0001000011011101", 25836 => "1000100111001010", 25837 => "1111101000010010", 25838 => "0101110101111110", 25839 => "1100110101111011", 25840 => "0110010100100011", 25841 => "0101110000100111", 25842 => "0011111111010111", 25843 => "1010011110011001", 25844 => "0100000110001100", 25845 => "0111110000000101", 25846 => "0011101011011000", 25847 => "1000111110101100", 25848 => "1100100100110101", 25849 => "1000111011110111", 25850 => "0110101100101101", 25851 => "0010010111011001", 25852 => "1000101100110101", 25853 => "0101110000101110", 25854 => "1111111111011100", 25855 => "0010100110111101", 25856 => "0111011010001101", 25857 => "0001111011000101", 25858 => "1111110010110001", 25859 => "1110101100001110", 25860 => "0010111110100100", 25861 => "0110010110100000", 25862 => "0010100001100010", 25863 => "1100010000110010", 25864 => "0010111101110101", 25865 => "1011011111100110", 25866 => "1001100010010000", 25867 => "1101010101000010", 25868 => "1010001001011011", 25869 => "0001111010100111", 25870 => "0000010001111011", 25871 => "0100001000110111", 25872 => "0000100000001011", 25873 => "0111001101010011", 25874 => "1000000011010000", 25875 => "1101101111011110", 25876 => "0010011111010011", 25877 => "0010010101001001", 25878 => "0001000001110110", 25879 => "0010001111000001", 25880 => "1101100011100100", 25881 => "0111010000001111", 25882 => "1100000001100110", 25883 => "1101100110001111", 25884 => "0111101000100000", 25885 => "1100011000011110", 25886 => "0111101101100101", 25887 => "0111000100010100", 25888 => "1110111010111100", 25889 => "1001010001010110", 25890 => "0011010110101000", 25891 => "0100110000110100", 25892 => "0001011111010110", 25893 => "1011001000101110", 25894 => "0000010100001110", 25895 => "0100010100001000", 25896 => "1100010111001100", 25897 => "1001111001011010", 25898 => "1010010011010101", 25899 => "0010011001101111", 25900 => "0010001100110001", 25901 => "0011100011111100", 25902 => "1111011001111011", 25903 => "0010000110111011", 25904 => "0111010011010001", 25905 => "1011010000001001", 25906 => "1011110100010011", 25907 => "1100001011000110", 25908 => "0100001100110000", 25909 => "0011011010010000", 25910 => "0011011111111011", 25911 => "0100000011000101", 25912 => "1111111000111110", 25913 => "1000000000110011", 25914 => "0111101111100101", 25915 => "0001000010101001", 25916 => "1001111000011001", 25917 => "1101111111000110", 25918 => "0100001010110010", 25919 => "1001110100011011", 25920 => "1010001010001001", 25921 => "0010110100101001", 25922 => "0010111111111011", 25923 => "1110100111000000", 25924 => "1011111101001111", 25925 => "1110110010101101", 25926 => "1011011011010011", 25927 => "1001010000110000", 25928 => "0101001101110001", 25929 => "0010011011111111", 25930 => "0000100010001000", 25931 => "0101111111011001", 25932 => "0111101000101110", 25933 => "0010111100110100", 25934 => "0100011000000011", 25935 => "1100101000010100", 25936 => "0111011011111110", 25937 => "0011111010011110", 25938 => "1110111100101110", 25939 => "0101010010101110", 25940 => "1000010111110111", 25941 => "1010011010110101", 25942 => "1110010011100011", 25943 => "1011011110010000", 25944 => "1001001111011101", 25945 => "1011010101101010", 25946 => "0000001010000010", 25947 => "0010111100000001", 25948 => "1000100101110011", 25949 => "0110111110111001", 25950 => "0011001011010010", 25951 => "0000011011111000", 25952 => "1100000011110101", 25953 => "0000000101100001", 25954 => "1101111110010011", 25955 => "0101101110101111", 25956 => "1011010001101011", 25957 => "0101110010100000", 25958 => "1101010010001100", 25959 => "1000101011111111", 25960 => "1011010010110100", 25961 => "0011010101010010", 25962 => "0000101111010010", 25963 => "1101000100100001", 25964 => "1110101101000110", 25965 => "1100000100100100", 25966 => "0111011110011011", 25967 => "0110001111001011", 25968 => "0000010010100010", 25969 => "1000111101011101", 25970 => "1111001011110101", 25971 => "1101101010010010", 25972 => "0101101001000110", 25973 => "0111001110110001", 25974 => "1110101011101000", 25975 => "1001001100001100", 25976 => "0101000110000010", 25977 => "1010111000100100", 25978 => "1000110101100101", 25979 => "0111100001111101", 25980 => "1000101100100111", 25981 => "0011011011111000", 25982 => "0111110010010000", 25983 => "0101000101100001", 25984 => "1111111001001011", 25985 => "0110001100001110", 25986 => "0100000001001000", 25987 => "1100010011000111", 25988 => "0101011010000001", 25989 => "0101001110111110", 25990 => "1110110010100011", 25991 => "1110101100001110", 25992 => "1000000011011010", 25993 => "1101010000100010", 25994 => "1100001101001111", 25995 => "0000000110101001", 25996 => "1110110000100001", 25997 => "1000000000011000", 25998 => "0111110110101010", 25999 => "0010010001000011", 26000 => "0011100001100001", 26001 => "1100100100000101", 26002 => "0000110110110111", 26003 => "0110110101000100", 26004 => "1101001111110111", 26005 => "0010111001011010", 26006 => "1010111011011010", 26007 => "1101100010100000", 26008 => "0100101011110111", 26009 => "0001010011110001", 26010 => "1111000100010101", 26011 => "1111101000110010", 26012 => "1111100111101100", 26013 => "0011010010010101", 26014 => "0110110000001101", 26015 => "0000101111101011", 26016 => "0110010010110111", 26017 => "1001001101100111", 26018 => "0000110110100110", 26019 => "1100000001111110", 26020 => "0110010101100000", 26021 => "1111000011101110", 26022 => "0000100111010011", 26023 => "0110110110010011", 26024 => "0001101100011000", 26025 => "0010000110001011", 26026 => "0110100111001111", 26027 => "0001000111111111", 26028 => "0110001011111011", 26029 => "1110001011111000", 26030 => "0110101101110010", 26031 => "1111001101000110", 26032 => "0110011000011010", 26033 => "1111100001101010", 26034 => "1010111111001011", 26035 => "1100001101000000", 26036 => "1010011010100101", 26037 => "1111100111110111", 26038 => "0001000111011000", 26039 => "0011011000010011", 26040 => "0000101100100001", 26041 => "0011111101011111", 26042 => "0101110100011001", 26043 => "1110010110000011", 26044 => "1101101011100010", 26045 => "0110011110110001", 26046 => "1001000011000011", 26047 => "0101111111110010", 26048 => "0110010001111010", 26049 => "1100101001011000", 26050 => "0100100101011010", 26051 => "0000101101111011", 26052 => "1101110101001000", 26053 => "1110110101110001", 26054 => "1100000000011101", 26055 => "1111111111101110", 26056 => "1010011110000100", 26057 => "1110010110010011", 26058 => "0101101000000110", 26059 => "0101101111101101", 26060 => "1011010111110010", 26061 => "0011100101001010", 26062 => "0101001001010111", 26063 => "0100010001100101", 26064 => "0000000011111111", 26065 => "1101001100100000", 26066 => "0001011010100010", 26067 => "1000001000000100", 26068 => "0101011010101110", 26069 => "1010101110110100", 26070 => "0001011010111101", 26071 => "1011011101100110", 26072 => "0010001101001110", 26073 => "1101110101100111", 26074 => "1101000100101100", 26075 => "1100101001010110", 26076 => "1010100100111001", 26077 => "0000100001000110", 26078 => "0010001000010000", 26079 => "0010111101011100", 26080 => "1000100011111001", 26081 => "0010111011111000", 26082 => "1000000100111011", 26083 => "0110000001011010", 26084 => "1111001100011100", 26085 => "0110010101000001", 26086 => "1111011010101001", 26087 => "1101001100101101", 26088 => "0101101010010010", 26089 => "0000101000100001", 26090 => "1100110101100010", 26091 => "1110111101001010", 26092 => "0010011111111010", 26093 => "0100010001110110", 26094 => "1010011010001001", 26095 => "1111111011110001", 26096 => "0000101000100001", 26097 => "1110001010110010", 26098 => "1000010010100101", 26099 => "1110011100110011", 26100 => "0111110001000010", 26101 => "0000001111001010", 26102 => "1110110010000101", 26103 => "0111000001001010", 26104 => "0111010000101000", 26105 => "1010000010100011", 26106 => "0010000010101101", 26107 => "1111011001111000", 26108 => "0100010000011010", 26109 => "0000010100010000", 26110 => "1001101010111111", 26111 => "0000101000000101", 26112 => "1100001010111010", 26113 => "0100110000010100", 26114 => "1101000000100110", 26115 => "1010110110001111", 26116 => "1010010110101011", 26117 => "1101010100101011", 26118 => "0000011011011010", 26119 => "1111010110001001", 26120 => "0000010101111010", 26121 => "0000010101111000", 26122 => "0010110100000100", 26123 => "0110011111110111", 26124 => "1111101101110101", 26125 => "1101001111100101", 26126 => "0110111011111000", 26127 => "1100010100001000", 26128 => "0100111110011111", 26129 => "1100001110010111", 26130 => "0111000100100110", 26131 => "1011010010110001", 26132 => "1111111010110000", 26133 => "0000001000110011", 26134 => "0001000001000101", 26135 => "1101010010001111", 26136 => "1011000101110101", 26137 => "0000101100101010", 26138 => "1111011010011101", 26139 => "0101100000101110", 26140 => "1011110011111100", 26141 => "1100100011101001", 26142 => "0011101000011100", 26143 => "1111101010000110", 26144 => "0101101110111100", 26145 => "0010000110110111", 26146 => "1011011110111001", 26147 => "0101100100011011", 26148 => "1110111100111000", 26149 => "1110001110001100", 26150 => "1111111100110100", 26151 => "1110011010100101", 26152 => "1000101010110111", 26153 => "0110011110001111", 26154 => "0000111110001110", 26155 => "0011101001011011", 26156 => "0110010001001100", 26157 => "0101000110111101", 26158 => "0100100101101110", 26159 => "0111101111011000", 26160 => "0101101001100010", 26161 => "0000000010111010", 26162 => "0100110010001111", 26163 => "1010101101111011", 26164 => "1011100100010010", 26165 => "0111000011000001", 26166 => "1101111010011111", 26167 => "1100110110101110", 26168 => "1101001001100010", 26169 => "1100011000000000", 26170 => "1010111001000001", 26171 => "1100111011000101", 26172 => "1101110011001011", 26173 => "1110011010011000", 26174 => "0100100000001101", 26175 => "1101100111110010", 26176 => "0101110011111111", 26177 => "0111011110111000", 26178 => "0010111010011111", 26179 => "0000000000001011", 26180 => "0110010011010000", 26181 => "1000000101110101", 26182 => "0001101000000111", 26183 => "0001100111100000", 26184 => "1101001101101110", 26185 => "1100100001101000", 26186 => "0101111111000000", 26187 => "0001010001111011", 26188 => "0110010011010110", 26189 => "1110101000001111", 26190 => "1001001110101110", 26191 => "0101100110101100", 26192 => "0011101100010111", 26193 => "1010010110111110", 26194 => "0110010110000011", 26195 => "1111100000011000", 26196 => "1100100111000101", 26197 => "0101111111101011", 26198 => "1111011000001100", 26199 => "1011101010100111", 26200 => "0111110111100101", 26201 => "0101101111111011", 26202 => "0111011000101101", 26203 => "1110101001011000", 26204 => "0111101001010011", 26205 => "1101000001101101", 26206 => "1101010000001100", 26207 => "1000011111100001", 26208 => "0111010011001110", 26209 => "0111101110010101", 26210 => "1001001001000100", 26211 => "1101011100000111", 26212 => "1011000011101100", 26213 => "0101011011011010", 26214 => "1001000010110110", 26215 => "1000100111101110", 26216 => "1011001110001110", 26217 => "1110100010110101", 26218 => "0111011110101010", 26219 => "0100001111001010", 26220 => "0001100000001011", 26221 => "0110010110011010", 26222 => "0011100010011011", 26223 => "1111011011110010", 26224 => "1000100111001111", 26225 => "0000101100000011", 26226 => "0111100111110110", 26227 => "1100001010000110", 26228 => "1010010101001000", 26229 => "0010010011110011", 26230 => "1010010010100000", 26231 => "0000000111101011", 26232 => "0000110001100001", 26233 => "1100010010110000", 26234 => "0110000001111010", 26235 => "0110111011101111", 26236 => "0101001111010010", 26237 => "0000001001001110", 26238 => "0111111000011011", 26239 => "0000100001011101", 26240 => "0001101101001110", 26241 => "0000100111100111", 26242 => "0000110000100000", 26243 => "0001010111101111", 26244 => "0000000000110010", 26245 => "0100011110010011", 26246 => "0000010110010001", 26247 => "0011110000100001", 26248 => "1010100110010000", 26249 => "1110011110100010", 26250 => "0100001001011011", 26251 => "1011111011000101", 26252 => "1111011010110101", 26253 => "0011001011000001", 26254 => "0110011010101011", 26255 => "1111101011010011", 26256 => "1111111100111000", 26257 => "1110111111110011", 26258 => "1111001101010000", 26259 => "1101100000010110", 26260 => "1111100001010011", 26261 => "0010100011110011", 26262 => "0110100101101000", 26263 => "1000100111110111", 26264 => "1110011010100101", 26265 => "0101011010001011", 26266 => "0000100100100110", 26267 => "0110100001110000", 26268 => "0011100001000001", 26269 => "1111001101110000", 26270 => "1010011101011100", 26271 => "0000001000111000", 26272 => "0011110001001100", 26273 => "1000001010101001", 26274 => "0000101010011110", 26275 => "1100111110010011", 26276 => "1010011110101011", 26277 => "1100000101000011", 26278 => "0001001110111000", 26279 => "0011011110001111", 26280 => "1110000001010100", 26281 => "0011011010001110", 26282 => "0110011001001010", 26283 => "1111011001110111", 26284 => "0000000011101111", 26285 => "1111010110100010", 26286 => "0111100100001010", 26287 => "1101111010010011", 26288 => "0011100110110001", 26289 => "1110101110111011", 26290 => "0100010011111011", 26291 => "1101111110100101", 26292 => "0001100011111110", 26293 => "1011110001011011", 26294 => "1011110101101001", 26295 => "0100011011010110", 26296 => "0000111000000100", 26297 => "0011101001111001", 26298 => "1111101111101111", 26299 => "1000100000111110", 26300 => "1001000001111011", 26301 => "1111010011110101", 26302 => "1110100010010010", 26303 => "0111000110100001", 26304 => "1000010111110011", 26305 => "1101011010001000", 26306 => "1001011111100011", 26307 => "1000110010100111", 26308 => "0010110100010100", 26309 => "0100001111001001", 26310 => "1011011010001001", 26311 => "1101101101100111", 26312 => "0011110000001101", 26313 => "0111110101111101", 26314 => "0101010001001100", 26315 => "0100101100101111", 26316 => "0101001000101011", 26317 => "0001010010100100", 26318 => "0010000100101011", 26319 => "1101100011000010", 26320 => "1000010110101110", 26321 => "0101100101100001", 26322 => "0000001101011110", 26323 => "0101100100011011", 26324 => "0000011101111001", 26325 => "1000110001111101", 26326 => "1000001110001000", 26327 => "1110000100111101", 26328 => "1001011111100011", 26329 => "0001101010001001", 26330 => "0101001010011111", 26331 => "1010011010110010", 26332 => "0010001110010011", 26333 => "1000100111011011", 26334 => "0000100011001011", 26335 => "1100010110011010", 26336 => "1101001011101001", 26337 => "0110000011010000", 26338 => "1101000111011000", 26339 => "1111001101001101", 26340 => "1001000011011011", 26341 => "0110100001110111", 26342 => "0001111011101111", 26343 => "0101010010101010", 26344 => "1000101101100111", 26345 => "1100010111111011", 26346 => "1000011110011001", 26347 => "1101000010101010", 26348 => "1100111001101010", 26349 => "0101100010101110", 26350 => "0101110000000001", 26351 => "1111110111010111", 26352 => "1010100010011001", 26353 => "0010111111010001", 26354 => "0111010011000100", 26355 => "1110010000011000", 26356 => "0101100000010011", 26357 => "0001110111010001", 26358 => "0001010111110111", 26359 => "0111001010000001", 26360 => "1101001111010010", 26361 => "1100110111101111", 26362 => "1101101000001101", 26363 => "1100101101001101", 26364 => "1101010011011111", 26365 => "1011010001000000", 26366 => "1011010001010010", 26367 => "1100010011111000", 26368 => "1101001010100011", 26369 => "0000001001100011", 26370 => "1011101101110000", 26371 => "0100110101111001", 26372 => "0011010001100111", 26373 => "1010101111001001", 26374 => "0010111000010110", 26375 => "1110100111011000", 26376 => "1010001010100000", 26377 => "1110000101100000", 26378 => "0100000100001101", 26379 => "0101101001000110", 26380 => "0011101001001011", 26381 => "0000010001000001", 26382 => "0001101110110111", 26383 => "1010000100100011", 26384 => "1010011111100100", 26385 => "1000011110101101", 26386 => "1011101101000000", 26387 => "1111011111010010", 26388 => "0101100110110011", 26389 => "1010111110011000", 26390 => "0000000010100011", 26391 => "0111100001010010", 26392 => "1011110001011101", 26393 => "0100000000111101", 26394 => "0001001101110011", 26395 => "0000000001110101", 26396 => "1001011011110011", 26397 => "1100111011011110", 26398 => "0111001001011010", 26399 => "0101110111101101", 26400 => "1011010110011101", 26401 => "1011110011110011", 26402 => "0001100100001101", 26403 => "0111111000001110", 26404 => "0001000111100110", 26405 => "1100000111010010", 26406 => "0010011011000110", 26407 => "0101000101110001", 26408 => "1011101001001000", 26409 => "0101100101100011", 26410 => "1000110101100101", 26411 => "1001011100011010", 26412 => "0010000010100101", 26413 => "1011111011001010", 26414 => "0000011110110110", 26415 => "1100111000101110", 26416 => "1101001011110100", 26417 => "0010110111000101", 26418 => "0101010111001100", 26419 => "1000010100111001", 26420 => "0001001011000101", 26421 => "0110100101101111", 26422 => "0000101110011010", 26423 => "0111000100001101", 26424 => "1001101110010101", 26425 => "1101101010011101", 26426 => "0011101010101010", 26427 => "1100101010010100", 26428 => "1111010010001010", 26429 => "1001101011001011", 26430 => "1100000001111100", 26431 => "1111010010100010", 26432 => "0111111011111101", 26433 => "1100001110101100", 26434 => "0000110000000101", 26435 => "0101001011001001", 26436 => "1011101011000010", 26437 => "1011011011010010", 26438 => "1011000001011001", 26439 => "0010000100010001", 26440 => "0101000111011101", 26441 => "1010110011010010", 26442 => "1001110101111001", 26443 => "1011001110111010", 26444 => "0101001111111110", 26445 => "1000111110000011", 26446 => "1001001100101001", 26447 => "1000100011100110", 26448 => "0111001110010100", 26449 => "1101010100101111", 26450 => "1100010111010010", 26451 => "0111100101010111", 26452 => "0001001010001011", 26453 => "0010001100001111", 26454 => "0100010000011001", 26455 => "1010011011111011", 26456 => "1110100010000101", 26457 => "0101111011101110", 26458 => "1100101000110001", 26459 => "1000011100100011", 26460 => "0000001100010101", 26461 => "1011000110000111", 26462 => "1011101101100101", 26463 => "0100001001111110", 26464 => "1011111010111001", 26465 => "0000111010000011", 26466 => "1001011100111000", 26467 => "0001010000011110", 26468 => "0001000101100000", 26469 => "0101100011001000", 26470 => "0010010101010011", 26471 => "1011010111000011", 26472 => "1100000100110100", 26473 => "0100010011001111", 26474 => "0110111001101011", 26475 => "1001111110111111", 26476 => "0101010110100011", 26477 => "0101110111101100", 26478 => "0100101110101111", 26479 => "1100001111000001", 26480 => "1001000000100101", 26481 => "1100000001110100", 26482 => "0000001001110011", 26483 => "1001010011111110", 26484 => "1111111110001011", 26485 => "0100011000010110", 26486 => "0101101111100011", 26487 => "1010010111010010", 26488 => "0011001011010000", 26489 => "1110000011111100", 26490 => "1101000101101100", 26491 => "1011100010010100", 26492 => "1001100001101011", 26493 => "1010001011110011", 26494 => "0010101010100110", 26495 => "0010001100110100", 26496 => "1100101110001111", 26497 => "1000011011001101", 26498 => "1001000100101101", 26499 => "1001001011111011", 26500 => "0000110010100000", 26501 => "1101011100110011", 26502 => "0100011001110100", 26503 => "1110101110111010", 26504 => "1001100100110000", 26505 => "0101000111100011", 26506 => "0110100110000011", 26507 => "1110000001100100", 26508 => "1110100111000101", 26509 => "0100101101001101", 26510 => "0010100000011101", 26511 => "0110010111000000", 26512 => "1001010000101100", 26513 => "0000110100110010", 26514 => "1101101110101010", 26515 => "1010000000111000", 26516 => "0101110000011110", 26517 => "1001011111000101", 26518 => "0111100101111110", 26519 => "0110111011011110", 26520 => "0000011011110110", 26521 => "1010010111000001", 26522 => "0100111010000111", 26523 => "1100110101010001", 26524 => "1011010101101011", 26525 => "0111101001100111", 26526 => "1110000010110110", 26527 => "1011010111000111", 26528 => "1100111100100100", 26529 => "1110011110010001", 26530 => "1000000101010001", 26531 => "1111111001100001", 26532 => "1010100011101111", 26533 => "0100010010111111", 26534 => "1011011011011111", 26535 => "1110101100110010", 26536 => "1011000101011001", 26537 => "1110000011111111", 26538 => "0000000100111110", 26539 => "0110010101010010", 26540 => "1101111010001101", 26541 => "1101010011011100", 26542 => "1101100001101111", 26543 => "1010111010110010", 26544 => "0100100001011101", 26545 => "1111010101111111", 26546 => "1111001100110100", 26547 => "1110010010100000", 26548 => "1000101101100001", 26549 => "0000000101100000", 26550 => "1001101011011100", 26551 => "0001111010111111", 26552 => "0111100101001001", 26553 => "0000000110100110", 26554 => "0110110101011011", 26555 => "0110110010011011", 26556 => "1111011010011110", 26557 => "0010010100111010", 26558 => "0011110111110100", 26559 => "1000000001001000", 26560 => "0111001100000101", 26561 => "1000111011000000", 26562 => "0011001110010110", 26563 => "1110110101010010", 26564 => "0101011001110001", 26565 => "1011101010101100", 26566 => "1100100110000001", 26567 => "1010101011111001", 26568 => "1011000000011100", 26569 => "1001000111011101", 26570 => "1011011111110011", 26571 => "1001000011010111", 26572 => "0111100110001111", 26573 => "0001001111110111", 26574 => "1100001111101011", 26575 => "0000100111111001", 26576 => "0011101001100001", 26577 => "0010011001010101", 26578 => "0100010011011011", 26579 => "0111101110100010", 26580 => "1011001011111011", 26581 => "0010101000100011", 26582 => "0010001000100011", 26583 => "1011001000111100", 26584 => "1000100100001011", 26585 => "0100100100010010", 26586 => "1111011001100100", 26587 => "1111010011100001", 26588 => "1101111101010100", 26589 => "1001001110100001", 26590 => "1110101001011100", 26591 => "1111001101101000", 26592 => "0100111111101101", 26593 => "1100000000111100", 26594 => "1011000001000000", 26595 => "1001100011000000", 26596 => "1000110111101011", 26597 => "1000110101011100", 26598 => "0010000111010111", 26599 => "0011000000011111", 26600 => "1000000011101011", 26601 => "1010111011011101", 26602 => "0010011001110111", 26603 => "1111101000000101", 26604 => "0100010011101101", 26605 => "0010011100001110", 26606 => "0010001001101010", 26607 => "0110000100100110", 26608 => "1101001011110010", 26609 => "1011100110111011", 26610 => "0101100110111101", 26611 => "0010011111011111", 26612 => "0011100011011011", 26613 => "1111010110010001", 26614 => "1001110000011101", 26615 => "1000011111011001", 26616 => "1011110100110101", 26617 => "1010001000000000", 26618 => "1010110000000001", 26619 => "0010110010011011", 26620 => "1111100110100011", 26621 => "1100001010110010", 26622 => "1011011011100101", 26623 => "0100011101101111", 26624 => "0101111011100111", 26625 => "1100111011111110", 26626 => "0010000110111111", 26627 => "0100001100100011", 26628 => "0111011011101101", 26629 => "1010001010000100", 26630 => "1011010100100111", 26631 => "1000110000001011", 26632 => "0011001000000100", 26633 => "1101011000111010", 26634 => "0010000100100110", 26635 => "0101001110100110", 26636 => "0110101101001111", 26637 => "1100010111101010", 26638 => "1101000001110111", 26639 => "1001001111101100", 26640 => "0110101100011100", 26641 => "1000001111010111", 26642 => "0101000000101011", 26643 => "0110011101001000", 26644 => "0101011001010000", 26645 => "0010011001001101", 26646 => "0111000110100010", 26647 => "0101111110110001", 26648 => "0100000101100010", 26649 => "1101001110010100", 26650 => "0001101011110101", 26651 => "0001010000000011", 26652 => "0011010101111100", 26653 => "0011011010001110", 26654 => "0100100111101000", 26655 => "1100000010000011", 26656 => "1101100101011000", 26657 => "1011100111001010", 26658 => "0110011010000110", 26659 => "0011110110010010", 26660 => "1000101110011100", 26661 => "1100101101011000", 26662 => "0011100010100110", 26663 => "0010110111100100", 26664 => "1111011110110001", 26665 => "0001101010101110", 26666 => "0001101110100100", 26667 => "1000110111111101", 26668 => "1010101010001101", 26669 => "1001000111010100", 26670 => "1101001100010101", 26671 => "0011101100000101", 26672 => "0111011010111011", 26673 => "1001000101011001", 26674 => "0000100110011111", 26675 => "0011000011000001", 26676 => "0110011111100110", 26677 => "1011000001001011", 26678 => "1000011101010011", 26679 => "0110011110000010", 26680 => "0011101000110001", 26681 => "1010110101001110", 26682 => "0100101001101011", 26683 => "0101000000100001", 26684 => "0100001110000010", 26685 => "0011011011101111", 26686 => "0101010010110100", 26687 => "1011011000111011", 26688 => "1110111001000010", 26689 => "1000101000101011", 26690 => "1101010101100000", 26691 => "1111101101000001", 26692 => "1111011011000111", 26693 => "1101011111100111", 26694 => "0010010101100011", 26695 => "1110111011111010", 26696 => "0011011101000001", 26697 => "0010010111001000", 26698 => "1111001101111001", 26699 => "0111101111100110", 26700 => "0100011000011001", 26701 => "1111010010111001", 26702 => "0001001011100100", 26703 => "0100000001000000", 26704 => "1110111000000001", 26705 => "1010110010010011", 26706 => "1110111000110011", 26707 => "1010110011010110", 26708 => "0100010110101010", 26709 => "1000101111000101", 26710 => "0010010000011110", 26711 => "0101000101011001", 26712 => "1111011011111110", 26713 => "1101111100100111", 26714 => "0010010011100001", 26715 => "1100011001111010", 26716 => "0001110001101111", 26717 => "0001100101010001", 26718 => "0110111000000011", 26719 => "0100010000100001", 26720 => "0100111010011101", 26721 => "0101110111110111", 26722 => "1100101000011011", 26723 => "0111000001101000", 26724 => "0011011101001011", 26725 => "1010010111111011", 26726 => "0000001011111000", 26727 => "1101000001000001", 26728 => "1001001001011101", 26729 => "0010111011111010", 26730 => "0011001010011110", 26731 => "0111111101000110", 26732 => "1111101000001010", 26733 => "1101010101111000", 26734 => "1000111100100011", 26735 => "0100101110111111", 26736 => "1011111011011011", 26737 => "0110010000111001", 26738 => "0100001101100011", 26739 => "0010100010100011", 26740 => "1101000011011011", 26741 => "1011000001000010", 26742 => "1011000111011100", 26743 => "1001111011100111", 26744 => "0111001010000111", 26745 => "0000011000100011", 26746 => "0001001011100001", 26747 => "1101001000010110", 26748 => "0000001100000010", 26749 => "1110011000110101", 26750 => "1111100110000001", 26751 => "0001000101001111", 26752 => "0011011101001000", 26753 => "0011111000010011", 26754 => "0101110100010010", 26755 => "0001011100000010", 26756 => "0100100011011101", 26757 => "1000000111101111", 26758 => "1011001101101110", 26759 => "0111101101111101", 26760 => "0000100101101010", 26761 => "0011010011110000", 26762 => "0011110101110011", 26763 => "0000111100001111", 26764 => "1001110000100001", 26765 => "0100110001101001", 26766 => "0011111101110111", 26767 => "1000010001111000", 26768 => "1100101101010100", 26769 => "1101111011101001", 26770 => "0001111100111101", 26771 => "0001010100001111", 26772 => "0110110000101011", 26773 => "0100101101101001", 26774 => "0110101110111011", 26775 => "0101000001010000", 26776 => "1110000001010011", 26777 => "1001001110000000", 26778 => "0000010010110101", 26779 => "0111011100010100", 26780 => "0111101011010011", 26781 => "0001110011111110", 26782 => "1000101000101111", 26783 => "0010011100101010", 26784 => "0011101111111001", 26785 => "0010011000011110", 26786 => "0111111101110010", 26787 => "0101011001111101", 26788 => "0010000011100000", 26789 => "1111001001111000", 26790 => "1111101011111000", 26791 => "1100101011101110", 26792 => "1000111110100111", 26793 => "1010101100100011", 26794 => "0101111000010000", 26795 => "0110101101100000", 26796 => "0111101000001110", 26797 => "1000011110001010", 26798 => "0001001101011001", 26799 => "0111001101011010", 26800 => "1100100100011010", 26801 => "0100001111011110", 26802 => "1000000101100110", 26803 => "0110010100100101", 26804 => "0001111011110011", 26805 => "0100110101111101", 26806 => "1100010111100001", 26807 => "0100100110100010", 26808 => "0111010110000001", 26809 => "1111111011101010", 26810 => "0000111100100111", 26811 => "1001100000000001", 26812 => "0011110000110110", 26813 => "1111000000100100", 26814 => "1000101000100011", 26815 => "1101001100001010", 26816 => "1100010010101101", 26817 => "0000011110010000", 26818 => "0011101111000111", 26819 => "1100000101111110", 26820 => "0101000111001001", 26821 => "1001011010110011", 26822 => "0010100110101101", 26823 => "0100110110111001", 26824 => "0100111011111110", 26825 => "0000110111000100", 26826 => "1100100100011110", 26827 => "0111011010010010", 26828 => "0111001101101101", 26829 => "0001010000110010", 26830 => "1111010010011110", 26831 => "1000010000010111", 26832 => "0011110001110110", 26833 => "0001101111010100", 26834 => "1010100110100001", 26835 => "0011110000001011", 26836 => "1000101101011000", 26837 => "1111000000001010", 26838 => "0000111111001101", 26839 => "0100101001111110", 26840 => "1111111111000110", 26841 => "1010010011100101", 26842 => "0011110100001011", 26843 => "1010010101011011", 26844 => "1001011110110010", 26845 => "1001100000100001", 26846 => "0100111011011101", 26847 => "0110001001010010", 26848 => "1001011001101110", 26849 => "0011111101110001", 26850 => "1001101010011110", 26851 => "1100100101001110", 26852 => "0110111110110111", 26853 => "0110110101001001", 26854 => "1000100010000111", 26855 => "1010111011011011", 26856 => "0111000101010110", 26857 => "1100000011111100", 26858 => "1100110111100111", 26859 => "1010101000100000", 26860 => "0111110000111101", 26861 => "1010111110110000", 26862 => "0010011110001110", 26863 => "1011110101000011", 26864 => "1110101100000111", 26865 => "1001111001010010", 26866 => "1010000011010010", 26867 => "1000001010110001", 26868 => "0000101000010101", 26869 => "1001100000100100", 26870 => "1110010111010101", 26871 => "1001011001011000", 26872 => "0101010011010101", 26873 => "1101001100111001", 26874 => "1110101011100001", 26875 => "0111010010010100", 26876 => "1100000100010111", 26877 => "0111110001110011", 26878 => "1101000100010111", 26879 => "0111010010101000", 26880 => "1100100010111111", 26881 => "1001001111010110", 26882 => "1111000000001010", 26883 => "0111000110110111", 26884 => "0001010010101110", 26885 => "1001110011101111", 26886 => "1010001110111010", 26887 => "0100101000000100", 26888 => "0101000001000101", 26889 => "1010001001111010", 26890 => "1101000000111110", 26891 => "0000011010010000", 26892 => "1001100101100011", 26893 => "1110111100111001", 26894 => "0011010001000111", 26895 => "1100010111111000", 26896 => "1100100100010101", 26897 => "1011011110001111", 26898 => "0101011110111000", 26899 => "0011111010011011", 26900 => "0001111111111110", 26901 => "1101110101101110", 26902 => "1010001110111000", 26903 => "0000010011000110", 26904 => "1110111101011100", 26905 => "0111111011111000", 26906 => "1100011010101010", 26907 => "1001110010001000", 26908 => "1101000010010100", 26909 => "0010001001101000", 26910 => "1010111000101010", 26911 => "0010101101000111", 26912 => "0011011111001101", 26913 => "1111010010101101", 26914 => "1011010010011111", 26915 => "0101110011010000", 26916 => "1111111001000110", 26917 => "1000110010110011", 26918 => "1010110011110100", 26919 => "0101101100101010", 26920 => "0110100111011001", 26921 => "1001111101101010", 26922 => "1010010111001101", 26923 => "1011100000111101", 26924 => "0101000111011111", 26925 => "1111111111001110", 26926 => "0101000000010100", 26927 => "0001111000101111", 26928 => "1000000000110101", 26929 => "1110000110010011", 26930 => "1000110110000010", 26931 => "0001010100100000", 26932 => "1110010110010010", 26933 => "0000100100100011", 26934 => "1001001010100110", 26935 => "0111100100111001", 26936 => "0111010001000000", 26937 => "0101010100111010", 26938 => "1000111101100100", 26939 => "1010000001100010", 26940 => "1100110100100101", 26941 => "0011110000010101", 26942 => "0001111010011011", 26943 => "1000100000001110", 26944 => "0110011000110010", 26945 => "1001110111100011", 26946 => "0101000010000010", 26947 => "1100101010101101", 26948 => "1111111001110011", 26949 => "1000001011111100", 26950 => "0101010100111111", 26951 => "1001111100101011", 26952 => "0100010111010100", 26953 => "0010000100011011", 26954 => "1100111010110101", 26955 => "0000111000110001", 26956 => "0101000111000000", 26957 => "1001000101010110", 26958 => "0010010001101011", 26959 => "0001101101101001", 26960 => "1000110000010011", 26961 => "1100110010100010", 26962 => "0111100010000011", 26963 => "0010111111110001", 26964 => "1110011000110100", 26965 => "1011110010111001", 26966 => "0001101001111110", 26967 => "1011011010001101", 26968 => "0011101101110101", 26969 => "1100001000000110", 26970 => "1111101100000101", 26971 => "1000111010010000", 26972 => "1111110101100010", 26973 => "0110000001000001", 26974 => "1011000001110001", 26975 => "0001011111001010", 26976 => "0110001000100001", 26977 => "0000110001101010", 26978 => "0010111011000111", 26979 => "1010111101110000", 26980 => "1100010000001100", 26981 => "1100011001011100", 26982 => "1000001010000011", 26983 => "1010100000011011", 26984 => "0000100111010001", 26985 => "0100100111000100", 26986 => "1111001010111000", 26987 => "0101011001011011", 26988 => "0011110101101111", 26989 => "1001011000111011", 26990 => "1001110101101111", 26991 => "1000111101111111", 26992 => "0101101111011010", 26993 => "1001110110010100", 26994 => "1100010000111101", 26995 => "1001110100111010", 26996 => "1011001100011010", 26997 => "1100111110101011", 26998 => "1100110010101010", 26999 => "1100100001001110", 27000 => "1001110000011000", 27001 => "0010010110011101", 27002 => "0100000111110110", 27003 => "1110111010011001", 27004 => "1000010011001000", 27005 => "1110101000011101", 27006 => "0100110011001101", 27007 => "1011001110001000", 27008 => "1001100010100111", 27009 => "0001011110011100", 27010 => "0101111110111001", 27011 => "1110110101011101", 27012 => "1000011111011101", 27013 => "0111100100110100", 27014 => "1000011011001001", 27015 => "0000100101011101", 27016 => "1001101111011110", 27017 => "0000000100101110", 27018 => "1100101111111110", 27019 => "0101111100010101", 27020 => "0110110111011011", 27021 => "0110100110001101", 27022 => "0000111001001010", 27023 => "1100001111000010", 27024 => "1000111111100110", 27025 => "1111101111001011", 27026 => "1001000111010011", 27027 => "0001011111010010", 27028 => "0101110110010111", 27029 => "0110110011010010", 27030 => "0110101100010010", 27031 => "1111000101111011", 27032 => "0010111110110110", 27033 => "0001000000011001", 27034 => "0000000100100101", 27035 => "0101001010010110", 27036 => "0010000111001000", 27037 => "0001101100101011", 27038 => "0011100100010101", 27039 => "0001111011101001", 27040 => "1111100010000101", 27041 => "1000111110100111", 27042 => "1100011100100010", 27043 => "1110110110001010", 27044 => "1111100000001011", 27045 => "0010111011101010", 27046 => "0001000110111111", 27047 => "0111000001111100", 27048 => "1100000110000001", 27049 => "1001000110101000", 27050 => "1100110100011001", 27051 => "1001001000001100", 27052 => "0000000110111100", 27053 => "0011001011110110", 27054 => "1011010100001000", 27055 => "0010000010111101", 27056 => "1010011001110100", 27057 => "1100110011111100", 27058 => "1101100011001000", 27059 => "0111111101001101", 27060 => "0101000010001001", 27061 => "0011100010101100", 27062 => "0001000111011000", 27063 => "1111101110110100", 27064 => "1110010001111110", 27065 => "0011100010111000", 27066 => "0000011011001011", 27067 => "1001100000100000", 27068 => "1010101000000010", 27069 => "1110001111010000", 27070 => "0110010000011011", 27071 => "0011010101011000", 27072 => "1000100011100100", 27073 => "0010011100100100", 27074 => "0011110011010000", 27075 => "1000110010011010", 27076 => "1110011011010011", 27077 => "0011101001011101", 27078 => "0000100100111001", 27079 => "1110100100111000", 27080 => "1101100101101101", 27081 => "1011101100110010", 27082 => "1001001101111000", 27083 => "1100011000100001", 27084 => "0110010001011000", 27085 => "1101011011100101", 27086 => "0011010101010010", 27087 => "0000011001000101", 27088 => "0110000011110001", 27089 => "1011101110001000", 27090 => "1111111111101110", 27091 => "1101110010010011", 27092 => "0110100000111011", 27093 => "1010000001011110", 27094 => "1111000101001110", 27095 => "0100000000001110", 27096 => "0101000001001011", 27097 => "1010111110110001", 27098 => "0000111101000001", 27099 => "0000000010001010", 27100 => "0010000100110000", 27101 => "1100010100000010", 27102 => "0110010101011100", 27103 => "0010110010001111", 27104 => "0100010000010011", 27105 => "1000101001001001", 27106 => "0100101101010101", 27107 => "1101101100000110", 27108 => "1011110111110010", 27109 => "0010100100100011", 27110 => "0000000001001100", 27111 => "1100000100110011", 27112 => "1111000111101000", 27113 => "0011111010101000", 27114 => "1010110111110100", 27115 => "0100001111111100", 27116 => "1110000010100011", 27117 => "0011011001011010", 27118 => "0111000101010101", 27119 => "0011011001100000", 27120 => "1111011110101000", 27121 => "0001110011100010", 27122 => "1000011101001101", 27123 => "1000000100111010", 27124 => "1111010101000101", 27125 => "0000000001010000", 27126 => "1000110010101101", 27127 => "0101100110111010", 27128 => "0101110111011000", 27129 => "1011110100100100", 27130 => "0001010011011000", 27131 => "1110010110010111", 27132 => "1001011001100111", 27133 => "0011100101110010", 27134 => "1011001010010110", 27135 => "0101111010000111", 27136 => "0101001110100111", 27137 => "1100010000000001", 27138 => "1000001001110011", 27139 => "1100011101101010", 27140 => "1010010100001000", 27141 => "1100111101011011", 27142 => "1111000000001110", 27143 => "1011110010010011", 27144 => "1001111110010001", 27145 => "0011100000101000", 27146 => "1000110110110100", 27147 => "1111010001111110", 27148 => "0111100100010000", 27149 => "0111011000100010", 27150 => "0101111111101000", 27151 => "0011100100100101", 27152 => "1110110000100101", 27153 => "1011001010010110", 27154 => "1000110011110101", 27155 => "1101100100000001", 27156 => "0110111101100101", 27157 => "1100011101100001", 27158 => "0110001110000010", 27159 => "1111110001101000", 27160 => "0100111001011100", 27161 => "0111001111010010", 27162 => "1100010111100111", 27163 => "1111001101110011", 27164 => "0100101011001100", 27165 => "1000001000010100", 27166 => "1001111101000010", 27167 => "0010010001001000", 27168 => "0100100010101101", 27169 => "0011001100010001", 27170 => "1111001111100110", 27171 => "1100110110110110", 27172 => "0111010110101100", 27173 => "1111001001010111", 27174 => "0000110001101001", 27175 => "0010101000110010", 27176 => "1011111110001001", 27177 => "0111001010010011", 27178 => "1111100001110111", 27179 => "1001101100101110", 27180 => "0010011101000000", 27181 => "0111010010101001", 27182 => "0101001010010000", 27183 => "0001110101101100", 27184 => "1101100000011111", 27185 => "1000011110111000", 27186 => "1000101101001111", 27187 => "0111011011100100", 27188 => "0110111001100110", 27189 => "0001100101010000", 27190 => "0011101101101000", 27191 => "1100000010011010", 27192 => "1110001111000111", 27193 => "0000100101000111", 27194 => "0110001111111011", 27195 => "0010010111101011", 27196 => "0100000001111110", 27197 => "1000101110110001", 27198 => "1000000010001101", 27199 => "0101001101101011", 27200 => "0100100100100110", 27201 => "0011110000010010", 27202 => "1111111111000000", 27203 => "0011110101001100", 27204 => "0001001101010001", 27205 => "1111011110001111", 27206 => "1111010100100000", 27207 => "1011110100001100", 27208 => "0101101011000110", 27209 => "1011011100011001", 27210 => "0101110101111111", 27211 => "0101111101100000", 27212 => "1010001010011010", 27213 => "0111001101111101", 27214 => "0001100110100011", 27215 => "1010001111101011", 27216 => "1001000111010101", 27217 => "1111111010001100", 27218 => "1000111111011100", 27219 => "0010100111001110", 27220 => "0111101101001100", 27221 => "1001101101111010", 27222 => "1011010100100101", 27223 => "0111000101111111", 27224 => "0111100100111110", 27225 => "1000011111100010", 27226 => "1000000110100010", 27227 => "0000001011111100", 27228 => "1010110000101111", 27229 => "1110100010100100", 27230 => "1000011111100010", 27231 => "0101000101011101", 27232 => "0111010100011001", 27233 => "0110001000101111", 27234 => "1110010100110011", 27235 => "1010100001100101", 27236 => "1011011000000110", 27237 => "0100001001011111", 27238 => "1110111011110111", 27239 => "1100101010110010", 27240 => "0010110101111001", 27241 => "1110101011100101", 27242 => "1111110011110100", 27243 => "0100010001011011", 27244 => "0011110111011000", 27245 => "0000011110110111", 27246 => "1011001111001111", 27247 => "0011101011101110", 27248 => "0101001101010001", 27249 => "0110110000100110", 27250 => "1010110100101011", 27251 => "1000110100000011", 27252 => "1101001110101101", 27253 => "1000011111101001", 27254 => "0010011010011001", 27255 => "0101110001000000", 27256 => "1011010110001100", 27257 => "0101100110001111", 27258 => "0011001110100101", 27259 => "0111111010100001", 27260 => "0110100000001010", 27261 => "0110110110110100", 27262 => "0111010101100111", 27263 => "1111101010110010", 27264 => "1111011001000000", 27265 => "1000001011001100", 27266 => "0111110110111101", 27267 => "0011000000111010", 27268 => "1001011100100001", 27269 => "0110100011001101", 27270 => "1000110110011100", 27271 => "0001011101110010", 27272 => "0101010011000101", 27273 => "1000111111001011", 27274 => "0001110101001111", 27275 => "1011110010000000", 27276 => "1011001010110011", 27277 => "1111110101110010", 27278 => "0111100101100110", 27279 => "1001101000101110", 27280 => "1101010101110110", 27281 => "0110100000100101", 27282 => "0001010011110001", 27283 => "1110101111001110", 27284 => "0001110101111010", 27285 => "1111010010100000", 27286 => "1010100001101010", 27287 => "0111011001110111", 27288 => "1011110100000100", 27289 => "0111000101000000", 27290 => "0110111001011010", 27291 => "1101100010110101", 27292 => "0000010110001100", 27293 => "1110100111100101", 27294 => "0111100001110000", 27295 => "1000000010001010", 27296 => "0100011001111101", 27297 => "1011010001110000", 27298 => "1111111111010010", 27299 => "1010101010001010", 27300 => "0111010110110000", 27301 => "0001001010001111", 27302 => "1010110101000111", 27303 => "1000110101101001", 27304 => "0101011001101110", 27305 => "0011110000011101", 27306 => "0101101010010011", 27307 => "1111001011110101", 27308 => "1110001011000111", 27309 => "0101110101000000", 27310 => "0101000110011111", 27311 => "1010100011010010", 27312 => "1111110011010000", 27313 => "1011001111000001", 27314 => "0000100101100001", 27315 => "0011001100100101", 27316 => "1111111011100110", 27317 => "0001100010111100", 27318 => "1011100010010110", 27319 => "1011001010010011", 27320 => "1111000010010101", 27321 => "1111111101000000", 27322 => "1101010101100000", 27323 => "0010011110011101", 27324 => "0001100100001000", 27325 => "1111000011111011", 27326 => "1111001010000100", 27327 => "1010111110111100", 27328 => "0101110010010010", 27329 => "0111110001110100", 27330 => "1010011101000011", 27331 => "0101001110101100", 27332 => "0001100010101110", 27333 => "0101000001111010", 27334 => "1111001100011000", 27335 => "1100001000001011", 27336 => "1111001000010000", 27337 => "1001100001011010", 27338 => "1110110111111110", 27339 => "1100111000001000", 27340 => "0010111110110010", 27341 => "1001101011000001", 27342 => "0110000001101110", 27343 => "1000110000101110", 27344 => "0100100001100011", 27345 => "1110000010111010", 27346 => "1010111010101010", 27347 => "0010101101001001", 27348 => "0110000011100100", 27349 => "0100111000111100", 27350 => "1111001000001001", 27351 => "0111101000101010", 27352 => "1000110000101011", 27353 => "1010010100001011", 27354 => "1001011001000101", 27355 => "0101110111010111", 27356 => "1011000010000011", 27357 => "1001110000111110", 27358 => "1000101110100100", 27359 => "0011011100010000", 27360 => "1011111011000001", 27361 => "0000111010110111", 27362 => "1011100010100110", 27363 => "0111011110111101", 27364 => "0001111100100110", 27365 => "0111011001100000", 27366 => "0011011000110111", 27367 => "0111101010111100", 27368 => "0010101101001000", 27369 => "1011000011100011", 27370 => "0011011001001110", 27371 => "1111001011001011", 27372 => "0111111110101110", 27373 => "0101101011010010", 27374 => "1111011110110010", 27375 => "0011111110010111", 27376 => "1100011000101010", 27377 => "0010011100100001", 27378 => "1000110101100011", 27379 => "1101001110000110", 27380 => "0000100101000011", 27381 => "0111010001010100", 27382 => "0001001000111010", 27383 => "1001100110001101", 27384 => "0110000101101011", 27385 => "1011101100100101", 27386 => "1010101011101001", 27387 => "1001101011111110", 27388 => "1001110010010111", 27389 => "1100101010111001", 27390 => "1111100010011110", 27391 => "0111011111011111", 27392 => "0011111101000110", 27393 => "1101110010001100", 27394 => "1111001010110011", 27395 => "1010101000111101", 27396 => "1010011000010010", 27397 => "0110100100100110", 27398 => "1010010011110101", 27399 => "0100111111100011", 27400 => "1001000000101100", 27401 => "0100111101000101", 27402 => "0011101110001001", 27403 => "0010000000010000", 27404 => "1011001101010010", 27405 => "1101001111011000", 27406 => "0000010100001110", 27407 => "0100110000100111", 27408 => "0011111000011011", 27409 => "0001100001101010", 27410 => "0010011101001101", 27411 => "0000111000101010", 27412 => "0001110000001101", 27413 => "1000001000111101", 27414 => "0101111101100010", 27415 => "0110101000110011", 27416 => "0010001010101111", 27417 => "1101001111100110", 27418 => "0011110110101001", 27419 => "1010010101001000", 27420 => "0110000010101111", 27421 => "1101101101010010", 27422 => "0000010001011100", 27423 => "1001110001011001", 27424 => "0000110111000110", 27425 => "0011010111111011", 27426 => "0000000100111101", 27427 => "1001001100110000", 27428 => "0111001110010010", 27429 => "0100010000000011", 27430 => "0001110111100000", 27431 => "0001101100001100", 27432 => "0101111010000101", 27433 => "1000100101111010", 27434 => "1011110110001001", 27435 => "1000011001100101", 27436 => "0001111110001101", 27437 => "1110000110010010", 27438 => "0000010100101101", 27439 => "1010011000010010", 27440 => "0000111100001011", 27441 => "0011001111010001", 27442 => "1110011100001110", 27443 => "0111001001111011", 27444 => "0110010101010010", 27445 => "1001010010110111", 27446 => "0101110001100100", 27447 => "0101111100110010", 27448 => "0010011111111011", 27449 => "0000000110100101", 27450 => "0011110100110101", 27451 => "1001100011010101", 27452 => "1100001110111100", 27453 => "1111111000101000", 27454 => "1100110000010011", 27455 => "1011011110000001", 27456 => "1010010010011001", 27457 => "1001010011011011", 27458 => "0111111110100100", 27459 => "0001100001110101", 27460 => "0101010011101101", 27461 => "1001101100101011", 27462 => "1110011001110100", 27463 => "1111100010100110", 27464 => "0001011110001101", 27465 => "1101011000110010", 27466 => "0001110101100000", 27467 => "1100000000011001", 27468 => "1001111110011010", 27469 => "1011000010110000", 27470 => "1011100100001110", 27471 => "0111101001001111", 27472 => "0010110100100111", 27473 => "1111110000111111", 27474 => "0100011110001000", 27475 => "1010100101110010", 27476 => "0010100111001110", 27477 => "0001010000101100", 27478 => "0010100100110101", 27479 => "1010101000011100", 27480 => "0001111100000011", 27481 => "0010111110100001", 27482 => "0110111001110000", 27483 => "1000110001001000", 27484 => "0100001011000011", 27485 => "0100011001001111", 27486 => "1111010100100100", 27487 => "0010101101001001", 27488 => "0001101000000000", 27489 => "0110011001010111", 27490 => "1111010001111100", 27491 => "1011010011100011", 27492 => "1011000101000110", 27493 => "0101111100001110", 27494 => "0101110001110010", 27495 => "0111100000000101", 27496 => "1011100101011000", 27497 => "1001000101111110", 27498 => "1011001010010101", 27499 => "0111000010010110", 27500 => "1000100010101001", 27501 => "0111101111000010", 27502 => "1001001110110000", 27503 => "0111001111110100", 27504 => "0001110111100000", 27505 => "0011111000010101", 27506 => "1010000100100001", 27507 => "0011101111000000", 27508 => "1101100001101110", 27509 => "0111110011011111", 27510 => "1010010111110010", 27511 => "0001110101100010", 27512 => "0010001001111100", 27513 => "0110010011000111", 27514 => "1000001110010100", 27515 => "1101110111100111", 27516 => "0100011110001011", 27517 => "1110000011010111", 27518 => "0111000001101110", 27519 => "0001010101100100", 27520 => "1010100001000101", 27521 => "0001010011010101", 27522 => "0000100111101010", 27523 => "0111110010011110", 27524 => "0011100100011001", 27525 => "1001011100111101", 27526 => "1101001111001010", 27527 => "1010110111111110", 27528 => "1111111101000101", 27529 => "1101110000011110", 27530 => "0010111010101000", 27531 => "0110110010100011", 27532 => "1011001110111000", 27533 => "0111110001110001", 27534 => "0110111101100101", 27535 => "0011110100001001", 27536 => "1011110110101101", 27537 => "1001111000111000", 27538 => "0101011100111100", 27539 => "0111000110101011", 27540 => "1011010000100000", 27541 => "0101101110001110", 27542 => "0110001001011010", 27543 => "1110010110011111", 27544 => "0000101010101001", 27545 => "0101111110001100", 27546 => "1100100110000111", 27547 => "0010100011010011", 27548 => "1111111001100010", 27549 => "0001000001010110", 27550 => "1011001011100100", 27551 => "0011000001001001", 27552 => "0110101111001100", 27553 => "1100100011111110", 27554 => "0011100100000001", 27555 => "0101110011010011", 27556 => "0110000010110111", 27557 => "1001011000010100", 27558 => "1011000000001000", 27559 => "1110000011111110", 27560 => "1101010011101101", 27561 => "0110000101101011", 27562 => "1111110001100100", 27563 => "1100011010110010", 27564 => "0000000100001110", 27565 => "1001011111100000", 27566 => "0101100000000110", 27567 => "0110101000110110", 27568 => "1101000000000110", 27569 => "0001001101001110", 27570 => "0101001110101111", 27571 => "1000100100011011", 27572 => "1110110001000001", 27573 => "0011110110010110", 27574 => "0100010011100000", 27575 => "0011100000111100", 27576 => "0011100110111101", 27577 => "0001011011101101", 27578 => "0101101000001000", 27579 => "0101110101101011", 27580 => "0101010011000100", 27581 => "1001011100010011", 27582 => "1111010100010001", 27583 => "0101011101010100", 27584 => "1110110011010100", 27585 => "1111110001101100", 27586 => "0100000101111011", 27587 => "0100101000110011", 27588 => "0000101100001101", 27589 => "0000100011011001", 27590 => "0011011101101110", 27591 => "1010111010011000", 27592 => "1000100011010011", 27593 => "0100101000001011", 27594 => "0101011011100100", 27595 => "0001001100101111", 27596 => "1001100101011101", 27597 => "0001000000010110", 27598 => "0111011010000000", 27599 => "1010000100011111", 27600 => "0110011010000010", 27601 => "0110011001011001", 27602 => "0110001000100100", 27603 => "0001001101000110", 27604 => "1001011110000100", 27605 => "1101101111110111", 27606 => "0110101000110100", 27607 => "1110111101011110", 27608 => "1000000001011011", 27609 => "1100010001110101", 27610 => "1110000000000001", 27611 => "0100001101100100", 27612 => "0000000110110110", 27613 => "1000000100110111", 27614 => "1000000010011100", 27615 => "1011011110000000", 27616 => "1100010010000110", 27617 => "0111000011100000", 27618 => "0101011111001101", 27619 => "0000111101011110", 27620 => "1101100011101011", 27621 => "1010110111000110", 27622 => "1100100011111000", 27623 => "0010001010110110", 27624 => "0111000101001001", 27625 => "0000011100111011", 27626 => "0110101101000110", 27627 => "1100001000101111", 27628 => "0000101101000111", 27629 => "0101100010100110", 27630 => "1000111011000010", 27631 => "0010111111011101", 27632 => "0011010110001101", 27633 => "0010011000001101", 27634 => "1111010110100110", 27635 => "0101010001011000", 27636 => "0000001001100010", 27637 => "0111010110001101", 27638 => "0100100011001001", 27639 => "0011000101001100", 27640 => "1100100011110010", 27641 => "1001100101111111", 27642 => "1111110011010000", 27643 => "0111011001111100", 27644 => "0000101111100010", 27645 => "1000100010110110", 27646 => "1101010111011001", 27647 => "1111111001001100", 27648 => "0011100001101001", 27649 => "0000101100001110", 27650 => "1111101000110011", 27651 => "1011100011101011", 27652 => "1010010001010111", 27653 => "0000101001001110", 27654 => "1000010000100010", 27655 => "1000001110000011", 27656 => "1110000011010101", 27657 => "1100001110101001", 27658 => "0011011011010110", 27659 => "0001100011011100", 27660 => "1001000010100011", 27661 => "1110010111001111", 27662 => "1001000110011100", 27663 => "0011101001101110", 27664 => "1000111001111011", 27665 => "1011101000110100", 27666 => "1010111000011011", 27667 => "1111111110001011", 27668 => "1001111001011010", 27669 => "1000011111010101", 27670 => "0010110110110000", 27671 => "1110101011000000", 27672 => "0100011101001100", 27673 => "0101010100110011", 27674 => "0101100010100000", 27675 => "1011000001100111", 27676 => "1011110011111100", 27677 => "0011101010001100", 27678 => "0100000111111011", 27679 => "1011110101011010", 27680 => "1101001001001110", 27681 => "1011100100100111", 27682 => "1100001111101011", 27683 => "0000010000001111", 27684 => "1101010000110101", 27685 => "1000101000000001", 27686 => "0111101010000100", 27687 => "0101010110001010", 27688 => "0000000111110110", 27689 => "1101000101110110", 27690 => "1001111100110000", 27691 => "0101100101001110", 27692 => "1010110101010100", 27693 => "1001101010011111", 27694 => "1111000111010011", 27695 => "0011010001100010", 27696 => "1111100111100010", 27697 => "0101100000011100", 27698 => "1001011111111011", 27699 => "0011100101110010", 27700 => "0010010111100101", 27701 => "1001110101110010", 27702 => "0110111001010001", 27703 => "1000110110011000", 27704 => "0110110011100110", 27705 => "0101111001100101", 27706 => "1110001001010000", 27707 => "0111111101101001", 27708 => "1011011011111100", 27709 => "1000111101010010", 27710 => "0000011100100001", 27711 => "1111111110110001", 27712 => "0101101011110011", 27713 => "1110111011000001", 27714 => "1110101100101100", 27715 => "0110011011100101", 27716 => "0001011100111110", 27717 => "1100010000001110", 27718 => "1111011111011100", 27719 => "0110111011010001", 27720 => "1100000110111010", 27721 => "0110111101010011", 27722 => "0100101011111111", 27723 => "0011010111011010", 27724 => "0011011001011101", 27725 => "0001011010011100", 27726 => "1111100000010011", 27727 => "1100101101110000", 27728 => "1101000001100001", 27729 => "0010101110101101", 27730 => "0001100000101101", 27731 => "0111011111010101", 27732 => "1010110000101010", 27733 => "0000010110101101", 27734 => "0100010011101101", 27735 => "1011010010000011", 27736 => "1111000110010100", 27737 => "1011010001010110", 27738 => "0011010111100110", 27739 => "1110100000001011", 27740 => "1110101100111001", 27741 => "0010110011010000", 27742 => "0110110010001110", 27743 => "0100010111110100", 27744 => "1000110111100001", 27745 => "0110011100000110", 27746 => "1000100010011100", 27747 => "0110011101100001", 27748 => "1101100001111010", 27749 => "1100010000101010", 27750 => "1101100110100010", 27751 => "0011010011101010", 27752 => "1111010101100001", 27753 => "1011111100100010", 27754 => "1110001101011001", 27755 => "0000100010110111", 27756 => "0000110010001111", 27757 => "0011010000110001", 27758 => "1101110111111001", 27759 => "1110111000011100", 27760 => "0111000011000100", 27761 => "1101110011110100", 27762 => "1010000000010110", 27763 => "0100011111100000", 27764 => "0000111001111010", 27765 => "0001000110101010", 27766 => "0101010111011100", 27767 => "0001000111101001", 27768 => "0001100001111100", 27769 => "0100111111110011", 27770 => "0000000111111101", 27771 => "0101100011000100", 27772 => "1101110100101010", 27773 => "0110011111100000", 27774 => "0110100111101010", 27775 => "1001000101101011", 27776 => "0101011100000110", 27777 => "0100110001101010", 27778 => "0000100111010000", 27779 => "0011000010011011", 27780 => "1000111010001000", 27781 => "0001011000000000", 27782 => "1100010001100111", 27783 => "0011110110010100", 27784 => "1100101000101100", 27785 => "0110111010101110", 27786 => "0000001100010101", 27787 => "1110010001001101", 27788 => "1010110011101011", 27789 => "1010010001010011", 27790 => "0000110111011000", 27791 => "0010000110101011", 27792 => "1110110010101101", 27793 => "0010110000100111", 27794 => "0011100011010001", 27795 => "1101000101001100", 27796 => "0111110111110001", 27797 => "1011010011111100", 27798 => "0010111000101111", 27799 => "1110000101101000", 27800 => "1010100111001010", 27801 => "0000100001111001", 27802 => "1111101001001000", 27803 => "0110100010110001", 27804 => "0001001011010110", 27805 => "0101101101100010", 27806 => "1100010011000101", 27807 => "1000100100100010", 27808 => "0100110100000101", 27809 => "0010110001110011", 27810 => "1100100011010010", 27811 => "1110000000111101", 27812 => "0001011011100000", 27813 => "1100001101001110", 27814 => "0010010111000111", 27815 => "1011010100111101", 27816 => "1010110111001101", 27817 => "0000110110110110", 27818 => "0010100111101111", 27819 => "1010000110000001", 27820 => "0010010110110010", 27821 => "1101000000011110", 27822 => "1101000010110010", 27823 => "0010110001000101", 27824 => "1010001110010100", 27825 => "0001111111111010", 27826 => "0111001010010110", 27827 => "1000010001001001", 27828 => "1110011100001110", 27829 => "1100000111011101", 27830 => "0101111001111010", 27831 => "0110101000000110", 27832 => "0000110111000011", 27833 => "1011011000111011", 27834 => "0110101000111011", 27835 => "1010000011101100", 27836 => "1001010001010000", 27837 => "1111000101011110", 27838 => "1001011110010100", 27839 => "1010110001110000", 27840 => "0110010001001001", 27841 => "0011100111011110", 27842 => "0100100110011010", 27843 => "1100001100110001", 27844 => "0101100100100001", 27845 => "0000010000010001", 27846 => "1011000101000100", 27847 => "0111010111110011", 27848 => "0001100101110010", 27849 => "1001000010010111", 27850 => "1100110101100010", 27851 => "1111000111001000", 27852 => "1000101101000000", 27853 => "1011101000011001", 27854 => "0000100100000110", 27855 => "1110001111001000", 27856 => "1111000100110000", 27857 => "0111101001111000", 27858 => "1011010001101101", 27859 => "0001010010101010", 27860 => "0101011001011100", 27861 => "0010110111010011", 27862 => "1000001100010101", 27863 => "1100101110111011", 27864 => "0000101101001011", 27865 => "0110011111111000", 27866 => "1001100010110010", 27867 => "1111010010000011", 27868 => "0000110010001001", 27869 => "0011100001100000", 27870 => "0100000001011110", 27871 => "0000010001101100", 27872 => "1010111100100101", 27873 => "1100001010000001", 27874 => "1010110101111001", 27875 => "0001010111110111", 27876 => "1101011101111011", 27877 => "1101111011110001", 27878 => "0010110011010001", 27879 => "0010001110001010", 27880 => "0001110111111011", 27881 => "0010111110000011", 27882 => "1011100110010010", 27883 => "1001010011011100", 27884 => "1010110110010110", 27885 => "0001010100110100", 27886 => "1011011110010101", 27887 => "0101010010011101", 27888 => "0000100110111010", 27889 => "0000111101111101", 27890 => "1110101011000100", 27891 => "0100111010001111", 27892 => "0000111011101010", 27893 => "1001000101101010", 27894 => "0101001100101110", 27895 => "1011110000101010", 27896 => "1101011011110101", 27897 => "0100011111101110", 27898 => "1111110010111000", 27899 => "0110011000010010", 27900 => "0100010111101111", 27901 => "1000001001010001", 27902 => "0100000001100000", 27903 => "0101100001000101", 27904 => "0010110010000000", 27905 => "1100001001100000", 27906 => "1001011011100000", 27907 => "0000000000101101", 27908 => "0001000010000111", 27909 => "1011000100100100", 27910 => "0000000011100010", 27911 => "0010100010100011", 27912 => "0110101010100000", 27913 => "0010000100100100", 27914 => "0110011001101100", 27915 => "0101001101100000", 27916 => "1011010001000101", 27917 => "1010010000100000", 27918 => "1110100100010010", 27919 => "1110111111000101", 27920 => "1111101100010011", 27921 => "1010001101110010", 27922 => "0011000110011101", 27923 => "0000000111101000", 27924 => "0010001110010001", 27925 => "0100100111110111", 27926 => "1110110010010001", 27927 => "1000110011010110", 27928 => "0011011110001011", 27929 => "0000011111101110", 27930 => "1000110010000111", 27931 => "0011001111011100", 27932 => "0101000011011110", 27933 => "0110011000010111", 27934 => "0010100001110110", 27935 => "0001000001011111", 27936 => "1100101110110101", 27937 => "1000011000110001", 27938 => "0101000101100111", 27939 => "0100100011011111", 27940 => "0001011110010101", 27941 => "0100010001111101", 27942 => "0110111010111000", 27943 => "1111001000100001", 27944 => "1100101010010100", 27945 => "1101100111001010", 27946 => "0110110110011100", 27947 => "1101111000101011", 27948 => "1010101011000110", 27949 => "1110000100001000", 27950 => "1101001111100001", 27951 => "1001110001010000", 27952 => "0100010100101001", 27953 => "1000110001100010", 27954 => "1100110001000111", 27955 => "1000000001010011", 27956 => "1111011010101110", 27957 => "0111001111010100", 27958 => "1101100100101111", 27959 => "1011011111101110", 27960 => "0110111011010000", 27961 => "0000100010100100", 27962 => "1101000000010000", 27963 => "1000000100010001", 27964 => "1010110111010110", 27965 => "1101001111010000", 27966 => "0000111100101100", 27967 => "0011001000001101", 27968 => "1111001000101010", 27969 => "1010110011001000", 27970 => "1111110101001001", 27971 => "0011011111110001", 27972 => "1010011001100111", 27973 => "0100110011111000", 27974 => "0111001111110001", 27975 => "0110101000110000", 27976 => "1111000001011110", 27977 => "0110000110011111", 27978 => "1110000000000010", 27979 => "1101110000101001", 27980 => "1001101000100000", 27981 => "1110101110111000", 27982 => "0110100011100001", 27983 => "1101101001010001", 27984 => "1011100111011110", 27985 => "1011101010011111", 27986 => "1000110110001110", 27987 => "0011100010001101", 27988 => "1101010011001111", 27989 => "1101111111001111", 27990 => "0000100111100110", 27991 => "1101011011111100", 27992 => "1000111111000011", 27993 => "0011011100010000", 27994 => "0011000111100011", 27995 => "0111010110010111", 27996 => "0001111111001110", 27997 => "0100111100111110", 27998 => "0011011011000100", 27999 => "0110100110101100", 28000 => "0000111111110111", 28001 => "1010001110100000", 28002 => "0100100111101100", 28003 => "0011101010010001", 28004 => "0011100001111111", 28005 => "1000011000011100", 28006 => "1110000011101110", 28007 => "0010100111100110", 28008 => "1011111000110001", 28009 => "1011011111100100", 28010 => "0011011100110001", 28011 => "0011100001100000", 28012 => "1011000101011010", 28013 => "1101001110000110", 28014 => "0010110000110101", 28015 => "1101000011010000", 28016 => "1101010001100111", 28017 => "1110010010101101", 28018 => "1010111011110110", 28019 => "1001111010011001", 28020 => "0010000001011110", 28021 => "0001101101110101", 28022 => "0111010101000011", 28023 => "0101001101101010", 28024 => "0011001000011011", 28025 => "0011010110010011", 28026 => "1110101010111011", 28027 => "1001011100001101", 28028 => "0001010111111111", 28029 => "0101111000000011", 28030 => "0001000011011010", 28031 => "0110100111110000", 28032 => "0011000010001110", 28033 => "1111000111001001", 28034 => "1001011101100100", 28035 => "0110000001010010", 28036 => "1100001001111001", 28037 => "1010101000100111", 28038 => "0010111101110111", 28039 => "1100110101000011", 28040 => "0011000101100001", 28041 => "1100010010111000", 28042 => "0110010011101000", 28043 => "1101101100010100", 28044 => "0001110010111111", 28045 => "1110110000101110", 28046 => "1101010100100110", 28047 => "0100110001001101", 28048 => "1011111100111101", 28049 => "0000100100111101", 28050 => "1110011011111111", 28051 => "0000111111101110", 28052 => "1000100111001001", 28053 => "1001110111011110", 28054 => "1111101101011000", 28055 => "1111011101110110", 28056 => "0101010100000011", 28057 => "1100100000000011", 28058 => "1000011011000111", 28059 => "1001111100001100", 28060 => "1100100000010010", 28061 => "0001001111100100", 28062 => "0010101111110110", 28063 => "1110110001001101", 28064 => "0100101001000101", 28065 => "0010001111101101", 28066 => "1101101000000110", 28067 => "0101110001101101", 28068 => "1000010110111111", 28069 => "1101011111001110", 28070 => "1101100000110110", 28071 => "1100010100101100", 28072 => "1110001100010010", 28073 => "1000011000100111", 28074 => "1011010110111000", 28075 => "1010011000100101", 28076 => "0111001110011111", 28077 => "0010100001011100", 28078 => "1001010101111000", 28079 => "1010000101001010", 28080 => "1001010110010100", 28081 => "0100111010001110", 28082 => "1010011110011101", 28083 => "1110101000010011", 28084 => "1001111001011000", 28085 => "0010001010100111", 28086 => "1101111000101010", 28087 => "0010100101010000", 28088 => "1010110111100000", 28089 => "0100100111011110", 28090 => "0000011111110001", 28091 => "0001010011010111", 28092 => "1100000011000011", 28093 => "1111011110100001", 28094 => "0111000011010001", 28095 => "0000010011101000", 28096 => "0100001110001000", 28097 => "0100101000100100", 28098 => "1001011111101011", 28099 => "0101110010111000", 28100 => "0110100101000000", 28101 => "0000010000111111", 28102 => "0011011101001001", 28103 => "0001111101001110", 28104 => "0111110101100010", 28105 => "1111010010100111", 28106 => "1111000100101001", 28107 => "0111110101111001", 28108 => "0111101111011100", 28109 => "1011000001000010", 28110 => "0010101111111001", 28111 => "1000011110110110", 28112 => "1001010111000010", 28113 => "0011011100000100", 28114 => "0100111001100011", 28115 => "0011111000001010", 28116 => "0001001000111000", 28117 => "0110101101010100", 28118 => "0110010011101001", 28119 => "1110011101101011", 28120 => "0101010010000011", 28121 => "1011011001000101", 28122 => "1001111100001011", 28123 => "0001111100100111", 28124 => "0011100111111000", 28125 => "1011110101111011", 28126 => "1000100010000100", 28127 => "0011100110110010", 28128 => "1000101010110100", 28129 => "1001110111011111", 28130 => "1101011001100110", 28131 => "1001100011000001", 28132 => "1010001010011010", 28133 => "1000000111010111", 28134 => "0111010011110010", 28135 => "0101011000111101", 28136 => "0010111001100001", 28137 => "1000100000011111", 28138 => "0000100001011001", 28139 => "0001100010110110", 28140 => "0111011011010011", 28141 => "1010101110010000", 28142 => "1101011111100001", 28143 => "1001000101110100", 28144 => "1011011110010001", 28145 => "1010110111111010", 28146 => "1010111101000010", 28147 => "1001110010010100", 28148 => "0001101000010100", 28149 => "0100101001110101", 28150 => "1010000011110110", 28151 => "0111100111001010", 28152 => "1111110001100110", 28153 => "1100010010001111", 28154 => "1010011101011000", 28155 => "1000011001011111", 28156 => "1001010111110011", 28157 => "1010111010101011", 28158 => "0010001000010011", 28159 => "1100101100111001", 28160 => "1110001101001100", 28161 => "0101001011101000", 28162 => "0110000110011011", 28163 => "1110010001010000", 28164 => "0000101001000110", 28165 => "0111100110111001", 28166 => "1111000011101111", 28167 => "0111001000100010", 28168 => "0010101110011011", 28169 => "0111010000001110", 28170 => "0111010111111110", 28171 => "1101000011010100", 28172 => "0101100110000011", 28173 => "1101001001111100", 28174 => "0001011001011011", 28175 => "0010111110100000", 28176 => "0011100100010100", 28177 => "1010011110000011", 28178 => "0111010011000011", 28179 => "1110110010000010", 28180 => "0010010100011010", 28181 => "0011110001000000", 28182 => "1001100011001010", 28183 => "1000110111110110", 28184 => "1110110010000111", 28185 => "0111101101110110", 28186 => "0101001110110101", 28187 => "0011011011101001", 28188 => "0011001111011101", 28189 => "0101011111111011", 28190 => "0001010101111100", 28191 => "0111111100001001", 28192 => "0110100110000010", 28193 => "1110010110010100", 28194 => "0100011001010010", 28195 => "1110110001110110", 28196 => "1100011010111111", 28197 => "1110001010110101", 28198 => "1110000001101011", 28199 => "0001001101110000", 28200 => "1101000001010001", 28201 => "1111110001000111", 28202 => "0010111001001101", 28203 => "0001110001011000", 28204 => "1011100011101101", 28205 => "1011001111100101", 28206 => "1010000001110110", 28207 => "0001100100111100", 28208 => "0100111000010111", 28209 => "0011001010010101", 28210 => "0110001001110000", 28211 => "1110010010000001", 28212 => "0111000000011110", 28213 => "1100110010111011", 28214 => "0110000110100001", 28215 => "1110010110101011", 28216 => "1101000000100101", 28217 => "1000011100011000", 28218 => "1101110100011111", 28219 => "0110101011011110", 28220 => "0010000101100010", 28221 => "1000101001110011", 28222 => "1011110111100100", 28223 => "0110000000110111", 28224 => "1110101101010111", 28225 => "0010100110110010", 28226 => "0010001011100110", 28227 => "0011110010111111", 28228 => "0010101000000011", 28229 => "1110100010000111", 28230 => "1110011110001101", 28231 => "1010010111000000", 28232 => "0001011011101010", 28233 => "0010100011011110", 28234 => "1001010010101110", 28235 => "1110101110001000", 28236 => "0001011111101100", 28237 => "0100010110111101", 28238 => "1110011110001001", 28239 => "0101101111101100", 28240 => "1000111100000101", 28241 => "0100100011111001", 28242 => "1001011110001000", 28243 => "0111010110101100", 28244 => "1101111100100001", 28245 => "1110011101010111", 28246 => "0010011110111001", 28247 => "1011101111000011", 28248 => "0100000100101110", 28249 => "1011001110011100", 28250 => "0101111111001010", 28251 => "1110110001000001", 28252 => "1000011101111011", 28253 => "0011111111010110", 28254 => "0000111100010110", 28255 => "1111011001001110", 28256 => "1011001100100100", 28257 => "0101010000110100", 28258 => "0101100110100010", 28259 => "0000000011111011", 28260 => "0110100100011010", 28261 => "1111100101111001", 28262 => "1010000101101100", 28263 => "1101001010000100", 28264 => "0011101110000011", 28265 => "0110011110111110", 28266 => "1110110110000001", 28267 => "1101110111100011", 28268 => "0001111100001111", 28269 => "1011101010000000", 28270 => "0111011111101110", 28271 => "1001110100010000", 28272 => "0011001010011000", 28273 => "0111000101001010", 28274 => "0001010000001111", 28275 => "0101111001101101", 28276 => "1111111010010101", 28277 => "0011110000000001", 28278 => "0011110010111101", 28279 => "0011000111110011", 28280 => "0011011011110100", 28281 => "1111001010011111", 28282 => "1000111111010111", 28283 => "1101010110111000", 28284 => "0011001011100001", 28285 => "0110101101101001", 28286 => "0000000010101001", 28287 => "0000001011000111", 28288 => "1010100000111110", 28289 => "1010010010000111", 28290 => "0101101101101001", 28291 => "0110001011001011", 28292 => "0100000010100111", 28293 => "0011100000011101", 28294 => "0100100010000110", 28295 => "0101100000011101", 28296 => "1101010111100001", 28297 => "0001111100111010", 28298 => "0001010010011000", 28299 => "1001000100100100", 28300 => "0010110110001001", 28301 => "1100110100011110", 28302 => "0100100101011100", 28303 => "1001110001010010", 28304 => "1100111111000010", 28305 => "1000000100010011", 28306 => "1101110100001100", 28307 => "1001111100110111", 28308 => "1001001111101101", 28309 => "1111100011101110", 28310 => "1001111001101011", 28311 => "1000001110110110", 28312 => "0001001110110111", 28313 => "1011111100110100", 28314 => "1101010100001111", 28315 => "0000010000000010", 28316 => "0110000010010001", 28317 => "1001111100111101", 28318 => "0001101111001111", 28319 => "1000001000110100", 28320 => "0000100111100010", 28321 => "1001011001000100", 28322 => "1101111111100100", 28323 => "0000101100001000", 28324 => "1101110111100000", 28325 => "1010101001100011", 28326 => "1111011010011110", 28327 => "0110001110111110", 28328 => "0000100011001101", 28329 => "1000101101101110", 28330 => "0001101000101101", 28331 => "1100111101011011", 28332 => "0110010011010011", 28333 => "0101111010001011", 28334 => "1111011001010111", 28335 => "1100100010010101", 28336 => "0111001011101101", 28337 => "0111100110001100", 28338 => "1000000000001001", 28339 => "1001010010001100", 28340 => "1011000000010110", 28341 => "1001111001001101", 28342 => "1101111100101101", 28343 => "1001000101011000", 28344 => "0000111011100000", 28345 => "1111011101101110", 28346 => "1110111101100110", 28347 => "0100000001000101", 28348 => "0000100000001111", 28349 => "0001100101000101", 28350 => "0000111111110001", 28351 => "1101101100001110", 28352 => "0101010010011111", 28353 => "1111001011101110", 28354 => "0011111010100010", 28355 => "0110101101110100", 28356 => "0100100000010100", 28357 => "0100000001011110", 28358 => "1110011111011011", 28359 => "0111100110100101", 28360 => "0010010100110011", 28361 => "0010110110001001", 28362 => "1010110000010000", 28363 => "1001111111110100", 28364 => "0010100000111000", 28365 => "0111110000010100", 28366 => "0100011001100001", 28367 => "0101111101110101", 28368 => "0110110011001000", 28369 => "0000011010010111", 28370 => "1000101011100100", 28371 => "0011000101001000", 28372 => "0110100100111001", 28373 => "0100010000011010", 28374 => "1000110010011000", 28375 => "1100001001011111", 28376 => "0011110110000011", 28377 => "0001100011111010", 28378 => "1100101010011011", 28379 => "1100010011101000", 28380 => "0011111001010001", 28381 => "1001100000101000", 28382 => "1100111101110111", 28383 => "1000100101011101", 28384 => "0001111110000101", 28385 => "1101101111001010", 28386 => "0011111010000100", 28387 => "1100110000010000", 28388 => "0101000100110000", 28389 => "1110110111101000", 28390 => "0001010001001110", 28391 => "1111001101001111", 28392 => "1100110011011001", 28393 => "1100110100111110", 28394 => "0110000101001110", 28395 => "1111101011111111", 28396 => "0011100110011000", 28397 => "1001000100111100", 28398 => "0001101110000101", 28399 => "1000001110011000", 28400 => "1011100000111000", 28401 => "0100111000010000", 28402 => "1001110001010010", 28403 => "1011010101111111", 28404 => "0101000000001111", 28405 => "1011111011110010", 28406 => "0110110001100101", 28407 => "1000111101001111", 28408 => "1101100000010101", 28409 => "1010101101111011", 28410 => "1000111011011000", 28411 => "0111011010011001", 28412 => "0111100001100101", 28413 => "1000111100010100", 28414 => "0100100000000011", 28415 => "1001011001001011", 28416 => "0000010100011101", 28417 => "1110101101101110", 28418 => "1110110011100000", 28419 => "0100110110010100", 28420 => "1011001011101000", 28421 => "0000110101001010", 28422 => "0110101010011010", 28423 => "0100100011000101", 28424 => "0111000010010011", 28425 => "0110010010101011", 28426 => "0111101000110011", 28427 => "0011010011000101", 28428 => "0011010010011100", 28429 => "1000111111111100", 28430 => "1111001111011010", 28431 => "1110101011101011", 28432 => "0111011000011101", 28433 => "1101101000001011", 28434 => "1011011010101111", 28435 => "1100110100101101", 28436 => "1011001101110000", 28437 => "0000100001101011", 28438 => "0111000010111111", 28439 => "1111000000011011", 28440 => "1011000100111111", 28441 => "1110111101010010", 28442 => "1001111000000010", 28443 => "0110001001100100", 28444 => "0100110010000100", 28445 => "1110100111001010", 28446 => "0011110111111011", 28447 => "0001011100011110", 28448 => "1100000010000101", 28449 => "0110010010110101", 28450 => "1101111100110001", 28451 => "0101111000100011", 28452 => "0000001101001101", 28453 => "1100110010111000", 28454 => "1101111101101101", 28455 => "0010100010000101", 28456 => "0111100000100101", 28457 => "1100110111100000", 28458 => "1000101011000110", 28459 => "0101010000111000", 28460 => "0001110001000000", 28461 => "0110000000001100", 28462 => "1100010001111111", 28463 => "1001111001011000", 28464 => "0011010010000101", 28465 => "0111000101101001", 28466 => "0011010000001000", 28467 => "0000101000000000", 28468 => "0111101001101001", 28469 => "0111000101010001", 28470 => "0001110010011011", 28471 => "0101111101101111", 28472 => "0010111100110000", 28473 => "1111111010001100", 28474 => "1011011101101010", 28475 => "1110111111000001", 28476 => "1010000101110100", 28477 => "1000010000100000", 28478 => "1100010101011111", 28479 => "1111000101101111", 28480 => "0001011011000010", 28481 => "1000110001010000", 28482 => "1100000010001101", 28483 => "0010110111000101", 28484 => "1001011111010100", 28485 => "0111011110000011", 28486 => "1000100101111010", 28487 => "0011000101100000", 28488 => "1001100001011101", 28489 => "0100111001110100", 28490 => "1010000010011010", 28491 => "1101111011010101", 28492 => "0110010110110000", 28493 => "0111110011001101", 28494 => "0011101100001101", 28495 => "1110000101010000", 28496 => "0111101100011000", 28497 => "1111011001111010", 28498 => "0001110111101100", 28499 => "1100111111100100", 28500 => "0111000111010001", 28501 => "0111000111010111", 28502 => "1101010001100110", 28503 => "0111111001111011", 28504 => "1100000111011010", 28505 => "0000111110101100", 28506 => "1101000010001001", 28507 => "1100111101100100", 28508 => "0100110101011000", 28509 => "0101011111001101", 28510 => "0011001000111100", 28511 => "0101101011110100", 28512 => "0010010111110100", 28513 => "0010000010001010", 28514 => "0000100011111010", 28515 => "1000010011010100", 28516 => "0111110100011010", 28517 => "1010010000101011", 28518 => "1001001100011111", 28519 => "1010001111101111", 28520 => "0011010100001001", 28521 => "0110001001000110", 28522 => "0101011000111100", 28523 => "1100101011100001", 28524 => "0111001100010000", 28525 => "0100000010100111", 28526 => "0101110001111111", 28527 => "1100101111100000", 28528 => "1101001110011001", 28529 => "0011010101011101", 28530 => "1101000000010011", 28531 => "0111100110100110", 28532 => "0111001110011111", 28533 => "1011110010111100", 28534 => "1110101010100000", 28535 => "0111110000010100", 28536 => "0011111101011000", 28537 => "1010011001101110", 28538 => "1111111110001111", 28539 => "1011000110000110", 28540 => "0011000101000101", 28541 => "1010110111010000", 28542 => "0101000101011101", 28543 => "0110000101101111", 28544 => "1101101011000001", 28545 => "0111000100110101", 28546 => "1111101111000001", 28547 => "0100100101011100", 28548 => "0000111001100011", 28549 => "0111011000011110", 28550 => "1111011100011010", 28551 => "1011011010001111", 28552 => "1110110100011110", 28553 => "1010100001110000", 28554 => "1000110000000010", 28555 => "0001111000110011", 28556 => "1001010100010111", 28557 => "1101001101011101", 28558 => "1001000000010010", 28559 => "0110101101001100", 28560 => "0100110111110001", 28561 => "0010101100011101", 28562 => "0111101101000111", 28563 => "1011001111101111", 28564 => "1000001100010001", 28565 => "1101001110001110", 28566 => "0010110101110010", 28567 => "1010111011000100", 28568 => "0100000000001011", 28569 => "1101010001001111", 28570 => "0100000000111111", 28571 => "1111101011110111", 28572 => "1101111100111110", 28573 => "1001001110000001", 28574 => "1101110011101100", 28575 => "0111111100010000", 28576 => "0100111100011000", 28577 => "1100101000100100", 28578 => "1010100101110110", 28579 => "1111111001011101", 28580 => "1110111100110000", 28581 => "0100000000011111", 28582 => "1000110101001100", 28583 => "0001111000111111", 28584 => "0000010011111001", 28585 => "1001001101101111", 28586 => "0110010000100101", 28587 => "0010001111011101", 28588 => "0001011001111011", 28589 => "1000001011000000", 28590 => "0101100001110101", 28591 => "0001011001011111", 28592 => "0110110111010110", 28593 => "1000000010001000", 28594 => "1101111111110110", 28595 => "0001001001111111", 28596 => "0000011010000100", 28597 => "1110101010101100", 28598 => "0100101110110010", 28599 => "1011111101011111", 28600 => "0100001100101101", 28601 => "1110000110011011", 28602 => "1110110010000000", 28603 => "0110000001110110", 28604 => "1111001001101000", 28605 => "1000110001110100", 28606 => "0100110111100011", 28607 => "1101110001001011", 28608 => "1011011001011011", 28609 => "0101001110111010", 28610 => "0001100010110110", 28611 => "1110010001001010", 28612 => "0011101011100110", 28613 => "0101001010001000", 28614 => "1111011010011011", 28615 => "1000001101101110", 28616 => "0001010110100011", 28617 => "1110111101011111", 28618 => "0111011110111010", 28619 => "0111100100111000", 28620 => "0000000000100110", 28621 => "1111010101000000", 28622 => "0101111000111000", 28623 => "0000100010010110", 28624 => "1001101101110010", 28625 => "1110100110000001", 28626 => "0001110010000011", 28627 => "0110110000100111", 28628 => "0000100100111001", 28629 => "1111100100100010", 28630 => "1010100101101000", 28631 => "0111100111101111", 28632 => "1000011110000111", 28633 => "0101001010010101", 28634 => "0111000100110001", 28635 => "0100011101001100", 28636 => "1010000111000011", 28637 => "0011000011001010", 28638 => "1110110110011001", 28639 => "0101100100101000", 28640 => "0011001001010000", 28641 => "1100000000100000", 28642 => "1001001011000011", 28643 => "1111000111000010", 28644 => "0101111011010000", 28645 => "1101100000010000", 28646 => "1110100010011001", 28647 => "0011110010011001", 28648 => "0111001011000110", 28649 => "1000000111001100", 28650 => "1110011101111110", 28651 => "0010111100010110", 28652 => "0010101110001001", 28653 => "0000001101100101", 28654 => "0100011111010011", 28655 => "0000101101000011", 28656 => "0000110101111011", 28657 => "0101101101111010", 28658 => "1111000001001100", 28659 => "0001101110001011", 28660 => "1101000010111000", 28661 => "0000001001111010", 28662 => "0110000110010010", 28663 => "0100100001111000", 28664 => "0100100000101110", 28665 => "1110111011111100", 28666 => "1101001101001010", 28667 => "0111100111000001", 28668 => "1110100010100111", 28669 => "1000001110110100", 28670 => "1110111100111011", 28671 => "1001001110100101", 28672 => "1111100011000011", 28673 => "0110000100010100", 28674 => "0001010011011110", 28675 => "1001111001011000", 28676 => "0100001110000011", 28677 => "0010100110010011", 28678 => "0001000011101010", 28679 => "0010110110000011", 28680 => "1100001100001100", 28681 => "1010100000100001", 28682 => "0101000101011101", 28683 => "0000000010100110", 28684 => "1001001011000101", 28685 => "0000101010011110", 28686 => "0010110011101011", 28687 => "0001011011011000", 28688 => "0000110111010110", 28689 => "1101010110000100", 28690 => "1011100101000110", 28691 => "0011110010000101", 28692 => "0011100111001011", 28693 => "0001111010000111", 28694 => "1110100101001111", 28695 => "0111100110011101", 28696 => "0001011111110011", 28697 => "1101010100000000", 28698 => "0010100001100011", 28699 => "1001111100000010", 28700 => "0101110010001101", 28701 => "0111101001100101", 28702 => "1100110110100101", 28703 => "1100110110001010", 28704 => "0101110010011100", 28705 => "0000100100101010", 28706 => "0011111000111100", 28707 => "1100100011110011", 28708 => "1100011111110010", 28709 => "1110101110100010", 28710 => "1111010000001011", 28711 => "0011100001001011", 28712 => "0110110001000001", 28713 => "0111001000111101", 28714 => "1111100000011000", 28715 => "1101000000011001", 28716 => "1100111001011000", 28717 => "1111010100000101", 28718 => "1000000001111010", 28719 => "0000000101110100", 28720 => "0111111010000000", 28721 => "0101111011111100", 28722 => "0101100011110100", 28723 => "0111111111101110", 28724 => "0000110111001111", 28725 => "0101001000110101", 28726 => "1100011010000001", 28727 => "1010011011110100", 28728 => "1101111101001010", 28729 => "1010001001011011", 28730 => "0111010011110001", 28731 => "0110101101001101", 28732 => "1111001100001011", 28733 => "1110000110001110", 28734 => "1100110111111011", 28735 => "1010110000110101", 28736 => "1111000011000010", 28737 => "0100110011011110", 28738 => "1101111101000100", 28739 => "1101101110110011", 28740 => "1101110010111110", 28741 => "0100000001101000", 28742 => "0110100001000111", 28743 => "1010010011100111", 28744 => "1101101010101001", 28745 => "1111111100101111", 28746 => "1111000110110000", 28747 => "1101110111001010", 28748 => "0001100101001101", 28749 => "0111011001000011", 28750 => "1110101110011001", 28751 => "1011110100101111", 28752 => "1110001110111111", 28753 => "0101000000011011", 28754 => "1111010000000111", 28755 => "1011100010111010", 28756 => "1110001010100001", 28757 => "0010110010000100", 28758 => "0111100111110111", 28759 => "0110010101000011", 28760 => "0011101100011111", 28761 => "0110000000110010", 28762 => "0011100111101010", 28763 => "0001101100001101", 28764 => "1111111100001001", 28765 => "1011101110011001", 28766 => "1010110100001000", 28767 => "0000011111000000", 28768 => "0011110001110110", 28769 => "1000101000100110", 28770 => "0101110010100011", 28771 => "0000110001100011", 28772 => "1100111000111000", 28773 => "0001100110111100", 28774 => "1101101000010100", 28775 => "0110011011000110", 28776 => "1011110100100011", 28777 => "1000011111101101", 28778 => "0101101010101111", 28779 => "0010110111111011", 28780 => "0101100011111110", 28781 => "1100110110110100", 28782 => "0001100100001001", 28783 => "1110010101000101", 28784 => "0000111000111110", 28785 => "0000011110001001", 28786 => "0110111111000011", 28787 => "0011000010101011", 28788 => "1111111011010011", 28789 => "0101111010010000", 28790 => "0000101111101101", 28791 => "1001101110001000", 28792 => "1101000100100100", 28793 => "0000000111100000", 28794 => "1010110100100110", 28795 => "1000101100000111", 28796 => "0001101001001110", 28797 => "1000101110100100", 28798 => "0100001011000011", 28799 => "0001111000101011", 28800 => "0000100000101110", 28801 => "0111111110011010", 28802 => "0101110110001001", 28803 => "0011110000010110", 28804 => "1100100101000011", 28805 => "1001011010011111", 28806 => "0111111001111011", 28807 => "1010101111110110", 28808 => "1010000101100010", 28809 => "0100001101111111", 28810 => "0010000001001010", 28811 => "0011011001000111", 28812 => "1110101001011001", 28813 => "1110101001110010", 28814 => "0000001011101010", 28815 => "0011000111000101", 28816 => "1001001011011110", 28817 => "1011111011010010", 28818 => "0010100100000011", 28819 => "1101110011011011", 28820 => "0000101100001110", 28821 => "0100111011111101", 28822 => "1011010101011100", 28823 => "1010101100110001", 28824 => "1100000010010110", 28825 => "1011011010011000", 28826 => "0110011101000100", 28827 => "1111111111101111", 28828 => "0111111101001010", 28829 => "0111111101110111", 28830 => "1110100010000111", 28831 => "0001111110000100", 28832 => "1101001011010010", 28833 => "1110000100101110", 28834 => "0000001001101111", 28835 => "1100111110110100", 28836 => "1100110100010110", 28837 => "0000100011000110", 28838 => "0111100010011101", 28839 => "1110111001110101", 28840 => "0001000101010010", 28841 => "0001000010000110", 28842 => "1001011101010001", 28843 => "1110010000100100", 28844 => "1011001010111110", 28845 => "1011001010001011", 28846 => "0100101111000000", 28847 => "0111011101001000", 28848 => "0000101000101100", 28849 => "0011111101100001", 28850 => "0100001011111010", 28851 => "0010111100111000", 28852 => "0101000010111011", 28853 => "0010010000010011", 28854 => "1010100000100010", 28855 => "1100000100001100", 28856 => "0001000110000110", 28857 => "1001110100001100", 28858 => "0110111110101010", 28859 => "1000101111100101", 28860 => "1101101000111011", 28861 => "0101001110110101", 28862 => "0110010101110101", 28863 => "1011001100101110", 28864 => "0101001101100101", 28865 => "1111101010010110", 28866 => "1101010111110101", 28867 => "1110000000101010", 28868 => "1100100000110011", 28869 => "1000001010110001", 28870 => "1111101010100010", 28871 => "0001100010011100", 28872 => "1000010011101000", 28873 => "1000111000101000", 28874 => "1001000111111100", 28875 => "0010110000101010", 28876 => "0001111101110111", 28877 => "0111011100010001", 28878 => "1101010010011111", 28879 => "0010001001101011", 28880 => "1101001111011101", 28881 => "1101000100000010", 28882 => "1101111000011010", 28883 => "0011001011000001", 28884 => "1110110001000110", 28885 => "0011011001111010", 28886 => "1001100111001111", 28887 => "0101111110001100", 28888 => "0011111000101000", 28889 => "0000000111001001", 28890 => "1111010100110110", 28891 => "1100010010011111", 28892 => "1011110111110110", 28893 => "1110100110110111", 28894 => "0000001000110011", 28895 => "1010010101100010", 28896 => "0110011010000110", 28897 => "1110000000011111", 28898 => "1010111000000101", 28899 => "0111110110110110", 28900 => "0001011011011111", 28901 => "0111000001010001", 28902 => "0100111011101100", 28903 => "1011010100011110", 28904 => "1000001000011110", 28905 => "0100000001111101", 28906 => "0101110110111000", 28907 => "0001001100101101", 28908 => "0010001100001011", 28909 => "1101000101111100", 28910 => "0111111111000100", 28911 => "1110111111001100", 28912 => "1111001000010101", 28913 => "1010101001101111", 28914 => "0110101000110010", 28915 => "1110000011010100", 28916 => "1010111110100011", 28917 => "1001010011110101", 28918 => "0010010111111101", 28919 => "1011100111010000", 28920 => "1110100110000011", 28921 => "1010010001011110", 28922 => "1010001111101111", 28923 => "1111111111001101", 28924 => "1111010100000111", 28925 => "0110111101101101", 28926 => "0100111101110110", 28927 => "0101110101100100", 28928 => "1001101011110101", 28929 => "0100011001001100", 28930 => "0011001111110010", 28931 => "0011001011100110", 28932 => "0010011000001110", 28933 => "1100011101001101", 28934 => "0110001101111001", 28935 => "0110110010011101", 28936 => "0011111001001001", 28937 => "0010010010101101", 28938 => "0010010011000011", 28939 => "1101110111100100", 28940 => "0010111000001101", 28941 => "1111110110110001", 28942 => "0010100010110110", 28943 => "0101010001111100", 28944 => "0011110110110110", 28945 => "1011011110101111", 28946 => "1000001010110001", 28947 => "1010011001101010", 28948 => "0011111101000101", 28949 => "1101101001100111", 28950 => "1110010011101110", 28951 => "1110011111011000", 28952 => "0100011011100001", 28953 => "0001100111100001", 28954 => "0101000100011100", 28955 => "0010001101011011", 28956 => "1010100110011110", 28957 => "1111100001001101", 28958 => "1101000110010011", 28959 => "0101111110111110", 28960 => "1001011110010111", 28961 => "1110001100011011", 28962 => "1100100011001011", 28963 => "0100110011011111", 28964 => "0110000001000001", 28965 => "1010101011001000", 28966 => "0100010110000000", 28967 => "1110000000011011", 28968 => "0001000011000111", 28969 => "1000101100110010", 28970 => "1110011000001001", 28971 => "1100000001101111", 28972 => "1111001111111011", 28973 => "1000001010111001", 28974 => "1011010000110000", 28975 => "0110101011011001", 28976 => "0001011111001011", 28977 => "0111010001100111", 28978 => "0011010010011111", 28979 => "0110000110100000", 28980 => "1001101010000100", 28981 => "1011000110011010", 28982 => "0000011000100010", 28983 => "0001010101001100", 28984 => "0101100100111010", 28985 => "1010101000011100", 28986 => "1011010011101001", 28987 => "0011000001111000", 28988 => "0011101010101100", 28989 => "0110011100111101", 28990 => "0001110110101000", 28991 => "0110101111011010", 28992 => "1011010010011101", 28993 => "0000010010011110", 28994 => "0011000011111100", 28995 => "1000101000000110", 28996 => "1011111110100100", 28997 => "0100001011011001", 28998 => "0110000000000011", 28999 => "0000110100011101", 29000 => "1110000110000010", 29001 => "0011000011110011", 29002 => "0100100001010010", 29003 => "1001011010101011", 29004 => "0100100101101011", 29005 => "1101111110001011", 29006 => "0001101110100010", 29007 => "0010000010011000", 29008 => "1110000101101000", 29009 => "0001101001010110", 29010 => "0110010010111000", 29011 => "0010010001000101", 29012 => "1111101001100110", 29013 => "0000111010010011", 29014 => "0101001001010011", 29015 => "1100110011000011", 29016 => "1110000101011100", 29017 => "0000000110011011", 29018 => "0101101010101011", 29019 => "1010111011001001", 29020 => "0010100011010101", 29021 => "1001000011111000", 29022 => "1001111001000100", 29023 => "0001110101100000", 29024 => "0111000011000001", 29025 => "0111000100101101", 29026 => "1000100110010110", 29027 => "1100110001011110", 29028 => "0101111000100001", 29029 => "1001010110011001", 29030 => "0010010100010101", 29031 => "0100011001110100", 29032 => "1000101010110000", 29033 => "0110111100001000", 29034 => "1000001011011110", 29035 => "0001101010100011", 29036 => "0011111100110110", 29037 => "1100001011011010", 29038 => "0101101010000010", 29039 => "1001110000101100", 29040 => "0100100001010001", 29041 => "0100000010101011", 29042 => "0100101110111100", 29043 => "1100011101001100", 29044 => "0011001010011011", 29045 => "0110100011011010", 29046 => "0101111001100101", 29047 => "1101101000001011", 29048 => "1101101111110011", 29049 => "1001110011011111", 29050 => "1001110110001111", 29051 => "1100010011111011", 29052 => "0101110111110101", 29053 => "0101110110001011", 29054 => "0100100010101001", 29055 => "0001001110001010", 29056 => "1101111100101101", 29057 => "1110001110111110", 29058 => "0100011110111011", 29059 => "1000101010010110", 29060 => "0111100111001001", 29061 => "0011111100101100", 29062 => "0101011011001001", 29063 => "1011110001000100", 29064 => "1110010010111001", 29065 => "1100111010111101", 29066 => "0011011001000111", 29067 => "1100010111001001", 29068 => "0101111111000101", 29069 => "0111110010010101", 29070 => "0111000000100100", 29071 => "1010100100010111", 29072 => "1101011010011111", 29073 => "0010100011011101", 29074 => "1101011001100010", 29075 => "0100110110111101", 29076 => "0101011100000010", 29077 => "1011001001101000", 29078 => "0010111110001100", 29079 => "0111001111111011", 29080 => "1011111110000110", 29081 => "0100101001010101", 29082 => "0011100010011100", 29083 => "0110011000011001", 29084 => "0000011100111101", 29085 => "0000001010111011", 29086 => "0000100001101111", 29087 => "0111110001001111", 29088 => "0101100110000100", 29089 => "0001001011010100", 29090 => "1011110010110001", 29091 => "0011111000001100", 29092 => "0110100100000100", 29093 => "1001010001101100", 29094 => "1111011101111011", 29095 => "1010010111000110", 29096 => "1000100010100011", 29097 => "1011111101001011", 29098 => "0010001100110010", 29099 => "1001100101101110", 29100 => "1111000100110010", 29101 => "0111110000110000", 29102 => "0100011110100001", 29103 => "1100111000011111", 29104 => "1101111100110000", 29105 => "0001001001100000", 29106 => "1011011111011010", 29107 => "1100011001101001", 29108 => "1111011001111101", 29109 => "0000011000011111", 29110 => "0011111000001110", 29111 => "1101101110001111", 29112 => "1101101110100010", 29113 => "1100110100100110", 29114 => "1011000101000111", 29115 => "1111001001100011", 29116 => "0110111111011110", 29117 => "1101101101111000", 29118 => "0111011100100001", 29119 => "0111111101001100", 29120 => "0000101000011110", 29121 => "0011110110101011", 29122 => "0000011000011010", 29123 => "1101011111000010", 29124 => "1111010010111011", 29125 => "0011000100010111", 29126 => "1001011011001101", 29127 => "0000110010010010", 29128 => "0101101000010010", 29129 => "0100111111100101", 29130 => "0100110001110011", 29131 => "1001010011101101", 29132 => "1111110011101000", 29133 => "1000100111101011", 29134 => "0101100011000001", 29135 => "0011011111010010", 29136 => "0110001010000111", 29137 => "1011010101011100", 29138 => "0000111110111111", 29139 => "0001100101100010", 29140 => "1000100010010110", 29141 => "1111100010001110", 29142 => "1101010010000110", 29143 => "0100111101101100", 29144 => "0101011111111110", 29145 => "1001100011001101", 29146 => "1111000111000111", 29147 => "0101101011111010", 29148 => "0001100101110010", 29149 => "0011111111110110", 29150 => "0000011110100111", 29151 => "0001000011111111", 29152 => "0000110101100000", 29153 => "0011001011111111", 29154 => "1010010110111111", 29155 => "1101000101000001", 29156 => "1000101110000000", 29157 => "1000110111110111", 29158 => "0101111101000011", 29159 => "0110011101011101", 29160 => "1101100111011001", 29161 => "0000101000101000", 29162 => "1110000000111010", 29163 => "1001010111100000", 29164 => "0000011001101010", 29165 => "0011000011101100", 29166 => "1010100110000000", 29167 => "1001000100011101", 29168 => "0000010110101001", 29169 => "0000011010011110", 29170 => "0111101110111001", 29171 => "1100010000100001", 29172 => "1101100000001100", 29173 => "1111101000000111", 29174 => "1010101111000010", 29175 => "0110011011001001", 29176 => "0010011110001101", 29177 => "1001111010000011", 29178 => "1111011011000111", 29179 => "0000110000110110", 29180 => "0110101000101000", 29181 => "1000101000001100", 29182 => "1010101001011110", 29183 => "1000110010111001", 29184 => "1100110000110010", 29185 => "0010000110110010", 29186 => "0111110011100010", 29187 => "1011101011000010", 29188 => "1001000001101010", 29189 => "0011100110100010", 29190 => "0100101110111101", 29191 => "1111001100011111", 29192 => "0010101100101110", 29193 => "1001101011001111", 29194 => "1101110011110000", 29195 => "0110001111101111", 29196 => "1101010001111100", 29197 => "0001110011101111", 29198 => "1110010011011101", 29199 => "0111000101101111", 29200 => "1110111111101011", 29201 => "0000010010111000", 29202 => "0110000011010000", 29203 => "1010011110111001", 29204 => "1001100111111001", 29205 => "0011011000001110", 29206 => "1101110111010111", 29207 => "0110111000100111", 29208 => "0001010001010101", 29209 => "1011010001010001", 29210 => "1001111001001100", 29211 => "0001000100101011", 29212 => "0001111010000010", 29213 => "1001010011011000", 29214 => "1110111001001011", 29215 => "0110010110010100", 29216 => "1000101111100000", 29217 => "1110001010011110", 29218 => "1100101100000111", 29219 => "0110001001110000", 29220 => "1110110000101101", 29221 => "1001010011011011", 29222 => "0101100000010010", 29223 => "0110110100111110", 29224 => "0000110001000000", 29225 => "0011000111011110", 29226 => "0110001101011000", 29227 => "1100110001101101", 29228 => "1110100111111011", 29229 => "1011100010111011", 29230 => "0101001010011111", 29231 => "0101100110011011", 29232 => "1000110011011100", 29233 => "0011011001111111", 29234 => "1011100000101101", 29235 => "1111111110100010", 29236 => "0110011011010110", 29237 => "1011001101010001", 29238 => "1110111101001010", 29239 => "1011100110110101", 29240 => "0101100000001011", 29241 => "0000001010011110", 29242 => "1011111101100111", 29243 => "0101010011100100", 29244 => "1011010001000101", 29245 => "1001111010110110", 29246 => "0010111111010011", 29247 => "1000110100101001", 29248 => "1001001111000100", 29249 => "0001111111011111", 29250 => "0001001110010011", 29251 => "1111101111101001", 29252 => "0010110111110100", 29253 => "1010010110101001", 29254 => "1011000010000111", 29255 => "0110110111001000", 29256 => "0000011100110010", 29257 => "1101111101011100", 29258 => "0001000100111111", 29259 => "0010100010110011", 29260 => "1101011001001001", 29261 => "0110001000011001", 29262 => "0100010111001101", 29263 => "1001000100011001", 29264 => "0100100100000000", 29265 => "1111100100010110", 29266 => "0100100110101010", 29267 => "1010001110101110", 29268 => "1010000100111011", 29269 => "1010101100100110", 29270 => "0001110111001100", 29271 => "1111001001100100", 29272 => "1000000000111101", 29273 => "1100101101100101", 29274 => "0101011111011111", 29275 => "0111011011101100", 29276 => "0001011000010111", 29277 => "1110000010110000", 29278 => "0011100100000110", 29279 => "1101000100010001", 29280 => "1001100111000001", 29281 => "1001000100010011", 29282 => "1000001011000100", 29283 => "0011100001100100", 29284 => "0101110110001011", 29285 => "0111101001100100", 29286 => "1011010000101010", 29287 => "0111100101110010", 29288 => "0010001100101010", 29289 => "0000001010101100", 29290 => "0111010010110011", 29291 => "1010110001010001", 29292 => "0000001101101101", 29293 => "0001001100101011", 29294 => "1000001010100100", 29295 => "0110100010110001", 29296 => "1101001101010100", 29297 => "1001101111100000", 29298 => "1101101010010100", 29299 => "1000011111110110", 29300 => "1111110000101011", 29301 => "0111000010110111", 29302 => "0011000011010010", 29303 => "1010111010011111", 29304 => "1101110001111101", 29305 => "0001110000001100", 29306 => "1100010001111000", 29307 => "0000110110110001", 29308 => "0100011011011001", 29309 => "1000001011001011", 29310 => "0111110110111110", 29311 => "1101110001011111", 29312 => "1000110110100101", 29313 => "0111001001010001", 29314 => "0000100011010101", 29315 => "1100111110110110", 29316 => "1100011011000001", 29317 => "1011111100100101", 29318 => "0100100101100101", 29319 => "0010000001111011", 29320 => "1010011100000100", 29321 => "0000010000001111", 29322 => "0011011011111011", 29323 => "1010011010100100", 29324 => "0010011001100111", 29325 => "1000100010010101", 29326 => "1111101000011011", 29327 => "0010100011011001", 29328 => "0111010000001010", 29329 => "0111100010101001", 29330 => "1000110100101010", 29331 => "1000010110101011", 29332 => "1101110010001101", 29333 => "0101001000001111", 29334 => "0101011000000111", 29335 => "1011011110101111", 29336 => "1011110001001110", 29337 => "1000011100001011", 29338 => "1000100010101011", 29339 => "1110000110101110", 29340 => "0011101010111010", 29341 => "0100001011100011", 29342 => "1100000000001111", 29343 => "1111010001100000", 29344 => "0010110110111101", 29345 => "0111110110011011", 29346 => "1011011111001011", 29347 => "1100101001110101", 29348 => "0111101001000011", 29349 => "1111010100011010", 29350 => "0011001011101011", 29351 => "1011001001000001", 29352 => "1110000110111101", 29353 => "0101010110111110", 29354 => "1111000110010111", 29355 => "0000100101011101", 29356 => "1011111100011100", 29357 => "1011111100111001", 29358 => "0101110110010111", 29359 => "1000001110111011", 29360 => "1011010101000101", 29361 => "1110110000101110", 29362 => "0011101100111011", 29363 => "0111000111100111", 29364 => "0010011001000001", 29365 => "0101011110111110", 29366 => "0101101100111000", 29367 => "1000011011111011", 29368 => "0011101001111010", 29369 => "0010110010011011", 29370 => "1101010100011101", 29371 => "1111100011011001", 29372 => "1110110110011100", 29373 => "0100011100001100", 29374 => "1000111001111110", 29375 => "1000011001000010", 29376 => "1000100010111101", 29377 => "1101111001000111", 29378 => "0010010110110100", 29379 => "0110110110110110", 29380 => "0011111101101110", 29381 => "0010010011101101", 29382 => "0010110001011101", 29383 => "0010001001001000", 29384 => "1001100011101010", 29385 => "0001101101111011", 29386 => "0110001010011111", 29387 => "0011110011110010", 29388 => "0001000110010101", 29389 => "1001100100111010", 29390 => "1100001111010011", 29391 => "0100001111101101", 29392 => "0100001011001010", 29393 => "1001001101001101", 29394 => "1110000010110010", 29395 => "0001010101000011", 29396 => "1000000001100001", 29397 => "0110111000011001", 29398 => "0010111111101011", 29399 => "1101010111000011", 29400 => "1011110110100001", 29401 => "1001011001101011", 29402 => "0001111110101110", 29403 => "1001101110011000", 29404 => "0000101110011100", 29405 => "0110101011101101", 29406 => "1110011110001000", 29407 => "0001000001011111", 29408 => "1000000010101000", 29409 => "1010111001001010", 29410 => "0000011100100010", 29411 => "0010110000111100", 29412 => "0001110001101010", 29413 => "1001110111010101", 29414 => "0000111110101000", 29415 => "0101000001000010", 29416 => "1000110010001001", 29417 => "1100000100111111", 29418 => "1000100010000011", 29419 => "1110011101000010", 29420 => "1011100110101001", 29421 => "1011110011111010", 29422 => "1111111010101100", 29423 => "1010101001100011", 29424 => "1100111000010110", 29425 => "0000010111000101", 29426 => "0010010111101110", 29427 => "0001001010010001", 29428 => "1111101101101001", 29429 => "0010011011011101", 29430 => "0000011001111110", 29431 => "1000010101010111", 29432 => "1001000000001101", 29433 => "0010101011101011", 29434 => "0010011100100011", 29435 => "1001111110110001", 29436 => "0100001011111011", 29437 => "1110110001011011", 29438 => "0100010111001110", 29439 => "0001011110100000", 29440 => "0010100011001100", 29441 => "0111000110111110", 29442 => "1010110010100000", 29443 => "1100100110111011", 29444 => "0011100001011011", 29445 => "1011000110100101", 29446 => "1011000000100110", 29447 => "1101100100110110", 29448 => "1011011100001011", 29449 => "1010101101000000", 29450 => "1001110000100010", 29451 => "1110010010000000", 29452 => "0111010000100101", 29453 => "0000011001011011", 29454 => "1111011101111010", 29455 => "0010001011001010", 29456 => "0001001011001110", 29457 => "0011000100101011", 29458 => "0110100010111111", 29459 => "0010001010000010", 29460 => "0011011010110111", 29461 => "1011111111110111", 29462 => "0100100100001011", 29463 => "0011101110111101", 29464 => "1011000101000111", 29465 => "0110101101100000", 29466 => "1101001111111100", 29467 => "1001001111001101", 29468 => "1101101011011011", 29469 => "1010110101010100", 29470 => "0001010010110001", 29471 => "1110100000011000", 29472 => "1101011111110011", 29473 => "0100010010000000", 29474 => "1001111001001011", 29475 => "1011011001110101", 29476 => "1110001111101110", 29477 => "0000001001101000", 29478 => "0011111101101011", 29479 => "0111000001100101", 29480 => "0110000100111001", 29481 => "0100101000001110", 29482 => "1101100001011011", 29483 => "0010111001100000", 29484 => "0001101011100001", 29485 => "0010010101000001", 29486 => "1001000111110001", 29487 => "0110000101101110", 29488 => "1100011111100100", 29489 => "1110011100101000", 29490 => "1111111101000010", 29491 => "0010001011001010", 29492 => "0101011101100010", 29493 => "0101110000110011", 29494 => "0111110011010010", 29495 => "1110111010101100", 29496 => "0000000000010010", 29497 => "1101111011010110", 29498 => "0010111010110011", 29499 => "1111111100010111", 29500 => "1101101110000110", 29501 => "1111000101010010", 29502 => "0101001011100000", 29503 => "0100011011111001", 29504 => "0100111000111100", 29505 => "0001111110001001", 29506 => "0101000011010010", 29507 => "0101001100110010", 29508 => "1001010110001001", 29509 => "1011000000101000", 29510 => "0011111010100010", 29511 => "1100010101000001", 29512 => "1110100001011011", 29513 => "0001111010110110", 29514 => "0010010100000011", 29515 => "1111000011110001", 29516 => "1011101011001100", 29517 => "0100010010101000", 29518 => "1001001100111000", 29519 => "1001100010000001", 29520 => "0100110111100110", 29521 => "1010111000010100", 29522 => "1010001110100001", 29523 => "0100111010001110", 29524 => "0111001010111010", 29525 => "1010110110110001", 29526 => "0110100001000010", 29527 => "0010011111100111", 29528 => "1111110000011001", 29529 => "1110100001100111", 29530 => "1010101011110001", 29531 => "0000010100000110", 29532 => "0000011011011010", 29533 => "0101011000111000", 29534 => "1010100100011110", 29535 => "0011100101110001", 29536 => "0001111000100100", 29537 => "1111110001101001", 29538 => "1111111110011011", 29539 => "0110110000110000", 29540 => "0001111111000001", 29541 => "1101011011111110", 29542 => "0111011111100111", 29543 => "1000110110110101", 29544 => "0110100001110101", 29545 => "1100111110101000", 29546 => "1010110110101100", 29547 => "1001010111011110", 29548 => "0110101110111100", 29549 => "1111111110111100", 29550 => "0100000010110001", 29551 => "1000001000011000", 29552 => "1101011000010000", 29553 => "1110000101111000", 29554 => "0110011000000101", 29555 => "1011110101101110", 29556 => "1111000011000101", 29557 => "1011100000110100", 29558 => "0101101111000001", 29559 => "0101011010111001", 29560 => "1010110011111000", 29561 => "1010011110101011", 29562 => "0100000001001001", 29563 => "0100010111101111", 29564 => "0101011001000110", 29565 => "0111101000001100", 29566 => "1101110101001100", 29567 => "1011100111011000", 29568 => "0110100000001110", 29569 => "1010011110100100", 29570 => "0110111011100011", 29571 => "1110000100011001", 29572 => "0101100010011000", 29573 => "1010011011001001", 29574 => "0000010101111010", 29575 => "0111001101100101", 29576 => "1111100000110011", 29577 => "0101010010000111", 29578 => "0000110111011111", 29579 => "1101000100001100", 29580 => "0000111111101010", 29581 => "0011000100110000", 29582 => "0000011100001001", 29583 => "1001100000100110", 29584 => "1010111000100100", 29585 => "1010100111111101", 29586 => "1001011111001010", 29587 => "1010110010011101", 29588 => "1100111110110100", 29589 => "0111100101110010", 29590 => "1010000011111100", 29591 => "0111001101001100", 29592 => "0101100101001001", 29593 => "0100000000000110", 29594 => "1100101001000001", 29595 => "1000101001010101", 29596 => "1010001110001000", 29597 => "1110010111101101", 29598 => "0011010110011101", 29599 => "1111101110000000", 29600 => "1110101100001000", 29601 => "1101111010010111", 29602 => "1101000100100110", 29603 => "0011111100110000", 29604 => "0000000010011110", 29605 => "0011001000111000", 29606 => "0100001001100110", 29607 => "1110111000011110", 29608 => "1100010111000000", 29609 => "0010010011000011", 29610 => "1110111011011110", 29611 => "0100011010011111", 29612 => "1100110011011100", 29613 => "0111001101010010", 29614 => "0011001000110110", 29615 => "0001100110111100", 29616 => "1111010001101111", 29617 => "1100100111110100", 29618 => "1111100011100100", 29619 => "1000010010001101", 29620 => "1000010111010100", 29621 => "1000001100000001", 29622 => "0101110101010111", 29623 => "1110000111000001", 29624 => "1011100110110011", 29625 => "1010111011111001", 29626 => "1101011010110111", 29627 => "0010110000011011", 29628 => "0111000011000001", 29629 => "0001101010001110", 29630 => "1110000000010101", 29631 => "1010000111001010", 29632 => "0011101100000011", 29633 => "1101001010011110", 29634 => "0110011010110111", 29635 => "0000101010011111", 29636 => "0001001111101100", 29637 => "0011010010100111", 29638 => "0000010001001001", 29639 => "0111100101010110", 29640 => "1101101001001110", 29641 => "1110011011001111", 29642 => "0111011100100010", 29643 => "0001110100000101", 29644 => "1111000011111101", 29645 => "1001110000000011", 29646 => "1111110000001101", 29647 => "1100000001100111", 29648 => "0111000110000001", 29649 => "0111101100111110", 29650 => "0110001010010110", 29651 => "1110100011101000", 29652 => "0000000001000110", 29653 => "1010011001011010", 29654 => "1010010101010011", 29655 => "0100100011000101", 29656 => "0011000000101110", 29657 => "0101101110001001", 29658 => "1011010010010111", 29659 => "0100011101000111", 29660 => "1010101110011011", 29661 => "0111100001000111", 29662 => "1110001111000000", 29663 => "0010110110001101", 29664 => "1101100000001011", 29665 => "1001110100110000", 29666 => "1100011000011010", 29667 => "1000001011101011", 29668 => "1111110100100101", 29669 => "0001101001011110", 29670 => "1111000110110100", 29671 => "0000101011101111", 29672 => "1011100101111010", 29673 => "0011100101001001", 29674 => "1111100011111011", 29675 => "0101011100000111", 29676 => "1101101100011111", 29677 => "1000011110110111", 29678 => "0000010010101010", 29679 => "0100010101001000", 29680 => "0010101000001100", 29681 => "0001000011101011", 29682 => "0011010100111000", 29683 => "1110011100101100", 29684 => "0001101101101000", 29685 => "0010100101110010", 29686 => "0111101111001100", 29687 => "1011111010010011", 29688 => "0111100011010011", 29689 => "0110111110010111", 29690 => "1111011010010000", 29691 => "1101111010101001", 29692 => "1111010111001100", 29693 => "1000101001100000", 29694 => "1001100000011100", 29695 => "0100101010000101", 29696 => "0100111000000101", 29697 => "1011001001011011", 29698 => "1101100010100110", 29699 => "1011001001001011", 29700 => "0111000110001000", 29701 => "1000011110011001", 29702 => "1110101101010001", 29703 => "1100111011101110", 29704 => "0011100111000101", 29705 => "1111000001100111", 29706 => "1001101100011110", 29707 => "0010010001001101", 29708 => "0111110101011101", 29709 => "1110101110110011", 29710 => "1100000110100011", 29711 => "1101001001001100", 29712 => "1101010100110100", 29713 => "0010101101101001", 29714 => "1000101000001011", 29715 => "1111011000010000", 29716 => "0011011111001000", 29717 => "1110001000001001", 29718 => "0010001110010010", 29719 => "0110011100010000", 29720 => "0010000000000001", 29721 => "1101011110111000", 29722 => "0101100001000011", 29723 => "1001000101101011", 29724 => "0100101000101011", 29725 => "0001101100001110", 29726 => "0010001011101101", 29727 => "0010011011110110", 29728 => "0001101011000100", 29729 => "0011111100101000", 29730 => "1001101111001010", 29731 => "1100110111000101", 29732 => "1001010010011000", 29733 => "1100100100010000", 29734 => "0100110100100011", 29735 => "0010011101100101", 29736 => "0010101010101001", 29737 => "0111011111011001", 29738 => "1001011100010101", 29739 => "0010010100100001", 29740 => "1001000100010111", 29741 => "0011010011111101", 29742 => "1111101110001101", 29743 => "1111010111001000", 29744 => "0000110101111110", 29745 => "0011011100101011", 29746 => "0011010010010001", 29747 => "1000011101000101", 29748 => "0100000011100000", 29749 => "0011010111011110", 29750 => "0011111011010001", 29751 => "0111100010001000", 29752 => "1110001101111110", 29753 => "0111100011000100", 29754 => "0111000101100100", 29755 => "0000111100011110", 29756 => "1010011001110011", 29757 => "1110101001100111", 29758 => "0111111010110000", 29759 => "1111110000010110", 29760 => "1110001011101001", 29761 => "1011011001101111", 29762 => "1110100000101001", 29763 => "1000011011011010", 29764 => "1110011000111001", 29765 => "1100011110100111", 29766 => "0001011100100101", 29767 => "0101011101000001", 29768 => "1101110100101101", 29769 => "0011001011110000", 29770 => "0000111101100001", 29771 => "1101010000110001", 29772 => "1011001111000000", 29773 => "1111110110001110", 29774 => "0011011110000001", 29775 => "1001001001001010", 29776 => "1100111001011001", 29777 => "1011000000110001", 29778 => "0110000000111001", 29779 => "1001101001000010", 29780 => "1001010001111000", 29781 => "0100010011001101", 29782 => "1001111100011101", 29783 => "0111100000000111", 29784 => "0000111001110101", 29785 => "1010001110101011", 29786 => "0101011011101110", 29787 => "1101101000111110", 29788 => "0001011100000010", 29789 => "1010011011100110", 29790 => "1100110010100010", 29791 => "0000001011001101", 29792 => "0100010100101011", 29793 => "0100001000100001", 29794 => "0010000010011011", 29795 => "0000111100001100", 29796 => "1110010101000110", 29797 => "1010101011110111", 29798 => "1010110110101100", 29799 => "0110000010001111", 29800 => "0110010101111110", 29801 => "0001011111000100", 29802 => "1100010110000101", 29803 => "1111001011110110", 29804 => "0000000111110010", 29805 => "1001000111010110", 29806 => "1111001101010100", 29807 => "1001010001010110", 29808 => "1001001011011111", 29809 => "0111010110000100", 29810 => "0001001100011110", 29811 => "0001000100000110", 29812 => "0001111111010000", 29813 => "0100100101101011", 29814 => "0110100001101001", 29815 => "1110101111011100", 29816 => "0101110110101011", 29817 => "1100011001000111", 29818 => "0110010010001011", 29819 => "1101111001100011", 29820 => "0111101101101000", 29821 => "0000000010010001", 29822 => "0101011000011110", 29823 => "1010001000101111", 29824 => "0111101111111111", 29825 => "1101101111010110", 29826 => "0011110111111000", 29827 => "1011111001110001", 29828 => "0010110010110010", 29829 => "1100000010111101", 29830 => "1110010011010010", 29831 => "1010010011011110", 29832 => "0101101111000010", 29833 => "1110100000101011", 29834 => "0100100111010001", 29835 => "1111111011101000", 29836 => "0001101111110001", 29837 => "0111110100000011", 29838 => "1000111000100110", 29839 => "0000010100101010", 29840 => "1010110111000110", 29841 => "0110000100101011", 29842 => "1010011010110100", 29843 => "0011001110110011", 29844 => "0111111001101101", 29845 => "1110111011110110", 29846 => "1111001111010000", 29847 => "1111011111101111", 29848 => "1111110111001010", 29849 => "0101101101010110", 29850 => "1110111000011010", 29851 => "0010101001001100", 29852 => "1111010011000100", 29853 => "0111100000110000", 29854 => "1011000101010000", 29855 => "0101101101011010", 29856 => "1010101010110100", 29857 => "1111000011000000", 29858 => "0000010011011101", 29859 => "1000101100111110", 29860 => "0101100001010000", 29861 => "1110001000101010", 29862 => "0111110000111110", 29863 => "1100000000010100", 29864 => "1010100011111101", 29865 => "1000110001001000", 29866 => "1010010110001010", 29867 => "1110110010010101", 29868 => "1000101000100100", 29869 => "1011011010010101", 29870 => "0100011100101001", 29871 => "1010101111000110", 29872 => "1111011001101101", 29873 => "1001000101101101", 29874 => "1000100101110001", 29875 => "0101100101101011", 29876 => "0101010100110111", 29877 => "1100001001111110", 29878 => "1011101001000101", 29879 => "0110100011000010", 29880 => "1111000010110100", 29881 => "0100000011111010", 29882 => "0000011110110101", 29883 => "1110100000010100", 29884 => "1011010011101101", 29885 => "1000010101101111", 29886 => "0101110111010111", 29887 => "1111101010101100", 29888 => "1000001001000010", 29889 => "0100110001001010", 29890 => "0110011001001100", 29891 => "0100111000010110", 29892 => "0100101110100110", 29893 => "0110100111001000", 29894 => "0100100110011101", 29895 => "0011011000101100", 29896 => "1001000101010110", 29897 => "1001011101000111", 29898 => "0110001111011001", 29899 => "1101011110101011", 29900 => "0001011100010110", 29901 => "0011000111000111", 29902 => "0101000110011001", 29903 => "1101001011111101", 29904 => "0010011011001110", 29905 => "1111101111010010", 29906 => "1011101111001101", 29907 => "1111111111001100", 29908 => "1101110000100001", 29909 => "1101001101011101", 29910 => "1000010011110110", 29911 => "1000010001011001", 29912 => "0110100101010000", 29913 => "1001001111100110", 29914 => "1101101010101000", 29915 => "1011010111000011", 29916 => "1101101110000111", 29917 => "0100101100111010", 29918 => "0001110001101100", 29919 => "1111000101111010", 29920 => "1110011101011111", 29921 => "0100111001111111", 29922 => "0011110110110010", 29923 => "1011010110010001", 29924 => "0101111110001100", 29925 => "1001011000111111", 29926 => "1100010011111110", 29927 => "0110001111000000", 29928 => "0110011001011101", 29929 => "0010010010000010", 29930 => "1100010100010101", 29931 => "1101011000101011", 29932 => "0011001101000100", 29933 => "1101011100011011", 29934 => "1010100101000011", 29935 => "1111011101001100", 29936 => "1010000101100011", 29937 => "1111001000011001", 29938 => "0001100101111010", 29939 => "0000011000100000", 29940 => "1010111100111011", 29941 => "0101000001101011", 29942 => "1100100100111111", 29943 => "1000100011100100", 29944 => "0100000101001101", 29945 => "0011000000111001", 29946 => "1111110111110001", 29947 => "1111100100000001", 29948 => "0010011000111000", 29949 => "1011010110101011", 29950 => "0110101010000100", 29951 => "0101111000011111", 29952 => "0001100011010011", 29953 => "0011100111001001", 29954 => "0101001000100001", 29955 => "1101111001000011", 29956 => "0110000010000110", 29957 => "0111111001010110", 29958 => "1011100101110000", 29959 => "0111010101100011", 29960 => "1011101000101100", 29961 => "1001111001110000", 29962 => "0111011101111001", 29963 => "1111011101110011", 29964 => "0001101001111000", 29965 => "1010010011000010", 29966 => "1010101011111011", 29967 => "1100010010011001", 29968 => "1000101000000011", 29969 => "1100010111111011", 29970 => "0111011010110100", 29971 => "0001010010000011", 29972 => "1111100110111001", 29973 => "1101101111010110", 29974 => "1011101010000100", 29975 => "1010010000110111", 29976 => "0111111101100100", 29977 => "0011110011111101", 29978 => "1010101111010111", 29979 => "0001111000000100", 29980 => "1111000010001100", 29981 => "0001010010010000", 29982 => "0011111001100101", 29983 => "0110000010100010", 29984 => "1001011010100000", 29985 => "1101100001110100", 29986 => "1000100001100111", 29987 => "1101111111110111", 29988 => "1010100010001010", 29989 => "0101001000011000", 29990 => "1110010010111001", 29991 => "0111101000011001", 29992 => "1101111110111100", 29993 => "0000000001001010", 29994 => "1001111111110100", 29995 => "1111000010111110", 29996 => "1000001111000100", 29997 => "0110001001101101", 29998 => "0110011101101010", 29999 => "0001111000000000", 30000 => "1101110010001110", 30001 => "1001101000100110", 30002 => "1011010010011101", 30003 => "1000110011010101", 30004 => "1000100000010111", 30005 => "0000011011100101", 30006 => "0010001001100101", 30007 => "1111101101011100", 30008 => "0001110000100011", 30009 => "0100100110000001", 30010 => "1001000011000010", 30011 => "1001110111001011", 30012 => "0110100000001000", 30013 => "0110000010111010", 30014 => "0000110101000000", 30015 => "1011111001100100", 30016 => "0101011010111100", 30017 => "1110011010100000", 30018 => "0011001000111000", 30019 => "0111010000001011", 30020 => "1110010011011000", 30021 => "1101010001011001", 30022 => "0010100101011111", 30023 => "1010111101110110", 30024 => "1111110100111000", 30025 => "1111101100000101", 30026 => "0011001100100100", 30027 => "1101010110110110", 30028 => "1000101001111101", 30029 => "0100100011111101", 30030 => "0001110110000101", 30031 => "0010101010010111", 30032 => "0111111001100101", 30033 => "0111000001110001", 30034 => "0001010110000110", 30035 => "0111011011101011", 30036 => "0101111101001101", 30037 => "0010000110111010", 30038 => "0000011011100111", 30039 => "0001111011001110", 30040 => "1111101010111001", 30041 => "1001101101100100", 30042 => "0111100001001001", 30043 => "0100111001000001", 30044 => "1011011100100001", 30045 => "1010011111110100", 30046 => "1101100101011011", 30047 => "1010110010111101", 30048 => "1111011100000001", 30049 => "1001101100110111", 30050 => "1101101010000000", 30051 => "0001100001100110", 30052 => "0101010001110010", 30053 => "1000000111101000", 30054 => "0111001111001011", 30055 => "0110001101001110", 30056 => "1000111010000000", 30057 => "1110101101011111", 30058 => "1110010011011111", 30059 => "1110111010101011", 30060 => "0101010100110101", 30061 => "1111001111110111", 30062 => "1011011000111001", 30063 => "1101011100011101", 30064 => "0111010001011110", 30065 => "0011100001001001", 30066 => "1100011101011000", 30067 => "1111110100111010", 30068 => "1001110010000011", 30069 => "0000000000101100", 30070 => "0101010000111101", 30071 => "1110010100111101", 30072 => "0101110100000101", 30073 => "1011110110100110", 30074 => "1010001011011100", 30075 => "0011111001101010", 30076 => "1101101101011100", 30077 => "0011100011011111", 30078 => "0111000110101101", 30079 => "0110110101000110", 30080 => "1001010110101010", 30081 => "1110000100010111", 30082 => "0010011100001101", 30083 => "0010011101100011", 30084 => "1010111001001101", 30085 => "0011110101001111", 30086 => "0111111000101001", 30087 => "1101010001101100", 30088 => "1100011101110000", 30089 => "0111110101100000", 30090 => "1100000100111000", 30091 => "0100101010001111", 30092 => "1010010010011010", 30093 => "0110111001101010", 30094 => "1101011100101000", 30095 => "1101011100110000", 30096 => "0111011111110000", 30097 => "0001100001110111", 30098 => "0101110001100111", 30099 => "1001101000100010", 30100 => "1000001010111011", 30101 => "0110100101111001", 30102 => "0111001010011100", 30103 => "1100110100010010", 30104 => "0100001111111010", 30105 => "0110111111110100", 30106 => "0010100100101011", 30107 => "0011110011110000", 30108 => "0110110100010000", 30109 => "1101010011011001", 30110 => "0111000001110001", 30111 => "0111000000111100", 30112 => "1011011110000001", 30113 => "1100101010101111", 30114 => "0000101100111000", 30115 => "0100111000100111", 30116 => "0101000110111011", 30117 => "1011111001110011", 30118 => "1011011000110010", 30119 => "0100001011100101", 30120 => "0101100000010111", 30121 => "0011010011011011", 30122 => "1000111011010000", 30123 => "0001011100010111", 30124 => "0110001111101100", 30125 => "0101110111100001", 30126 => "1110000100111010", 30127 => "0111100001100110", 30128 => "1101010100110100", 30129 => "1000100010100000", 30130 => "1000110101111110", 30131 => "1011101011101101", 30132 => "0111010110101000", 30133 => "1100000111010111", 30134 => "0000000010001100", 30135 => "0010010101010110", 30136 => "1001111011011111", 30137 => "0010010101010100", 30138 => "1011110101010000", 30139 => "1100101101011110", 30140 => "1011101011000011", 30141 => "0101110111111000", 30142 => "0110111110110111", 30143 => "1001000110111111", 30144 => "1100110011011000", 30145 => "1000110101010110", 30146 => "1001101111100101", 30147 => "1101110111110100", 30148 => "0100000101011101", 30149 => "0001011001100100", 30150 => "0010011111101010", 30151 => "0001000000100000", 30152 => "0110001100001010", 30153 => "0111111110011010", 30154 => "0110111000111101", 30155 => "0010011001111110", 30156 => "1001000100010101", 30157 => "0011001101100001", 30158 => "0110011111100010", 30159 => "1101101111000001", 30160 => "0111101010110011", 30161 => "1101001111111011", 30162 => "1111111111010111", 30163 => "1010101010110111", 30164 => "1011111110101101", 30165 => "1111000110101000", 30166 => "1001011010100001", 30167 => "0100011110001011", 30168 => "1100001001100111", 30169 => "1001011011011100", 30170 => "0010011111011101", 30171 => "0100000001011000", 30172 => "0110100011010000", 30173 => "0010000011100110", 30174 => "1111100000110101", 30175 => "0001010000011011", 30176 => "0011001100101000", 30177 => "1111101101000011", 30178 => "1010010010111000", 30179 => "0110011011001101", 30180 => "1010110001101011", 30181 => "0110110110011110", 30182 => "1101011110100111", 30183 => "1010100010110101", 30184 => "0010110111001001", 30185 => "0100111011001010", 30186 => "0110010000000101", 30187 => "0111010101011110", 30188 => "1001000100110001", 30189 => "0111101011101000", 30190 => "0110101101011100", 30191 => "0010110110101010", 30192 => "1010111110100110", 30193 => "0111110110101010", 30194 => "0011000011000001", 30195 => "1010111100100001", 30196 => "0100001110010000", 30197 => "0101011101110110", 30198 => "1001110101101100", 30199 => "1101101001011000", 30200 => "1001011111111111", 30201 => "0110101111001101", 30202 => "0111011100111100", 30203 => "1001110100010100", 30204 => "0001001011011100", 30205 => "0110000101000111", 30206 => "1001011010001010", 30207 => "1111110000110110", 30208 => "1010101001000110", 30209 => "0110101101001110", 30210 => "0011100111111111", 30211 => "1100001100111001", 30212 => "0001110000001011", 30213 => "0010000111011101", 30214 => "0010100011011001", 30215 => "1000000010100011", 30216 => "0111100111110010", 30217 => "0111110000000110", 30218 => "0110101000001110", 30219 => "0100110011010101", 30220 => "1101101110110011", 30221 => "1100010110011010", 30222 => "0101011111100010", 30223 => "0101111011001011", 30224 => "1101011001101111", 30225 => "0101001110111011", 30226 => "0010010000010110", 30227 => "0100101000101011", 30228 => "0111011111001110", 30229 => "1001000011010011", 30230 => "0101001101101110", 30231 => "1001000000100111", 30232 => "1010101110111000", 30233 => "0001001010111100", 30234 => "1000101111101011", 30235 => "1011000101100100", 30236 => "0111000111101110", 30237 => "0000010111010000", 30238 => "1010010111100001", 30239 => "1011110011111110", 30240 => "1110100011011100", 30241 => "1101001100100010", 30242 => "1010101000111010", 30243 => "0011001111010110", 30244 => "1111111000000100", 30245 => "0110100111010100", 30246 => "0011010100000100", 30247 => "1010111101110001", 30248 => "1000011111001100", 30249 => "0011001110101100", 30250 => "0100101010001001", 30251 => "0011011001010101", 30252 => "0100011100100010", 30253 => "0010111000011100", 30254 => "1001010000011100", 30255 => "0001100110101101", 30256 => "1011011001001001", 30257 => "0000110100000101", 30258 => "1110101111110010", 30259 => "0101101000101100", 30260 => "0011110011100110", 30261 => "0000100000110111", 30262 => "1001011010101010", 30263 => "0010101110011110", 30264 => "0010101011100101", 30265 => "0000100010100100", 30266 => "0101110001111010", 30267 => "1101110000110100", 30268 => "1010101000100100", 30269 => "0011111101001100", 30270 => "1011010001111011", 30271 => "1100000010100000", 30272 => "1100111011111001", 30273 => "0101010000011100", 30274 => "0110011000010011", 30275 => "1100000000000110", 30276 => "0100110011011110", 30277 => "0100111000010010", 30278 => "0001100001100110", 30279 => "0000010010000100", 30280 => "1100000001000010", 30281 => "0001101100011011", 30282 => "0010101011011110", 30283 => "1100110101000101", 30284 => "0110000101010111", 30285 => "1001110100110111", 30286 => "0100100000111100", 30287 => "0110101100011001", 30288 => "0010111111110001", 30289 => "0010100110100100", 30290 => "1000000111111001", 30291 => "1100011001110100", 30292 => "0010101100000101", 30293 => "0110111011110100", 30294 => "0100010101111111", 30295 => "0111010100010001", 30296 => "1100000000100100", 30297 => "0111001100000011", 30298 => "0110010100000100", 30299 => "1110100101001110", 30300 => "0110010111001111", 30301 => "1110101100101000", 30302 => "0101001001111110", 30303 => "1000111101100111", 30304 => "1100101111100000", 30305 => "1101101100000111", 30306 => "0110111011101111", 30307 => "1111001001010110", 30308 => "1010101110111101", 30309 => "0100010110110000", 30310 => "1010001011111111", 30311 => "1000010111100011", 30312 => "1000100010010111", 30313 => "1100001000111100", 30314 => "0000101111100101", 30315 => "1001011101110000", 30316 => "1010011101101101", 30317 => "0001010010001111", 30318 => "1011100000111101", 30319 => "1010000101001100", 30320 => "1110111100101111", 30321 => "1010111011011010", 30322 => "1111110111110101", 30323 => "1011000100000110", 30324 => "0010111001111001", 30325 => "0010100000110010", 30326 => "0110010111110111", 30327 => "0000110111000100", 30328 => "1010010010110011", 30329 => "1100101000000011", 30330 => "1110000110110110", 30331 => "1101110110100000", 30332 => "1100011110111001", 30333 => "1111110001000111", 30334 => "0001110100000011", 30335 => "0110000110011101", 30336 => "0101001111111001", 30337 => "0100100010010000", 30338 => "1100001000010000", 30339 => "0011101000110011", 30340 => "0101101010001111", 30341 => "0000010010010011", 30342 => "0001001000110000", 30343 => "0010111000010100", 30344 => "1010100101010100", 30345 => "0101100101110001", 30346 => "1011111011010010", 30347 => "1100000001101010", 30348 => "0001110010010001", 30349 => "1100010110110000", 30350 => "1010111011100100", 30351 => "1110110000101100", 30352 => "0001111010111101", 30353 => "1101010111011111", 30354 => "0110101010100000", 30355 => "0111000010000010", 30356 => "0101100010110001", 30357 => "1010101001011101", 30358 => "0111111111101101", 30359 => "0000111101101111", 30360 => "1101100101101110", 30361 => "1101010110000000", 30362 => "0010101001110110", 30363 => "1111110011001011", 30364 => "1111010100001000", 30365 => "0110000100011001", 30366 => "1000000011110010", 30367 => "0010011000011110", 30368 => "1100010111110011", 30369 => "1101001011001000", 30370 => "1101001001110110", 30371 => "0010110110110100", 30372 => "0101100001110011", 30373 => "1001101100111010", 30374 => "1110110110101111", 30375 => "0000010011000101", 30376 => "1111111000110100", 30377 => "0000101110111110", 30378 => "1100110101000110", 30379 => "0000100010111011", 30380 => "1011100111110010", 30381 => "1011100011101001", 30382 => "0000011010111111", 30383 => "1110011110101001", 30384 => "1000000101101011", 30385 => "0011111000101111", 30386 => "1000111011101011", 30387 => "0011000000001000", 30388 => "1001001100111000", 30389 => "1010011000111100", 30390 => "1100000001000101", 30391 => "1110010010100001", 30392 => "1111000101110100", 30393 => "0101001111010101", 30394 => "1100011111110001", 30395 => "1110011110011111", 30396 => "1110100001101000", 30397 => "1110000101111010", 30398 => "1111100001100101", 30399 => "0000110111011111", 30400 => "0010001010011010", 30401 => "0010110111001001", 30402 => "0001111110000111", 30403 => "1011101001100000", 30404 => "1110110010110101", 30405 => "1010011110000001", 30406 => "0010111001011100", 30407 => "0100111011001010", 30408 => "1110011111010001", 30409 => "1101100011000100", 30410 => "0011000011010101", 30411 => "0100110010110101", 30412 => "1000110010110000", 30413 => "1010111111011001", 30414 => "1101111010111111", 30415 => "1100010100110101", 30416 => "1000100011000100", 30417 => "0001111101010001", 30418 => "1111111111010000", 30419 => "0001111101001001", 30420 => "0110000010111001", 30421 => "0111100111011111", 30422 => "0111011010011000", 30423 => "1111101010011100", 30424 => "1101101010010100", 30425 => "0110011001010011", 30426 => "0000001101111111", 30427 => "1001101101101101", 30428 => "0111011011000001", 30429 => "0110110110100110", 30430 => "0111110100011111", 30431 => "0100010101110111", 30432 => "0010001010001111", 30433 => "1010000001001111", 30434 => "1110100100111100", 30435 => "1000110110010110", 30436 => "1110010101000011", 30437 => "1110101010110111", 30438 => "0100010001110001", 30439 => "0110001100000110", 30440 => "0100110011001110", 30441 => "0001000111111000", 30442 => "0010111101101000", 30443 => "0001000001010011", 30444 => "0111011111100110", 30445 => "0101110011000000", 30446 => "0111101100000111", 30447 => "1101001110100100", 30448 => "1101111100101100", 30449 => "1001011001010111", 30450 => "0001001010100011", 30451 => "0010101101110010", 30452 => "1100111100000110", 30453 => "0100101000100001", 30454 => "1010100000100111", 30455 => "0000110100011001", 30456 => "1001000011100100", 30457 => "1001110010001111", 30458 => "1000011111110111", 30459 => "0011011001001010", 30460 => "0100100101010110", 30461 => "0110100110011010", 30462 => "0110001111110101", 30463 => "1001100101110100", 30464 => "1000100001001010", 30465 => "0111100011101001", 30466 => "0101011011010000", 30467 => "0010010111011010", 30468 => "1100100111111011", 30469 => "0000101111100111", 30470 => "1010100111111011", 30471 => "1010100110001101", 30472 => "0101101001001000", 30473 => "0111000011101111", 30474 => "0100111110111010", 30475 => "1100010000000010", 30476 => "1111100000100111", 30477 => "0111011001000100", 30478 => "1000111101110011", 30479 => "0011100011000110", 30480 => "0101011101001110", 30481 => "0000110101110101", 30482 => "0010001001010001", 30483 => "0010111011010110", 30484 => "1010010110101001", 30485 => "0010100111000101", 30486 => "1000011011111000", 30487 => "1100010110110000", 30488 => "1011110100010100", 30489 => "0000110100001001", 30490 => "0001010011100101", 30491 => "1111001101111001", 30492 => "0010010101010100", 30493 => "1000110010101110", 30494 => "1001001111111100", 30495 => "1100001010101101", 30496 => "1101010100100100", 30497 => "1010011101001111", 30498 => "0101100011111101", 30499 => "1000100010101110", 30500 => "1000101111011011", 30501 => "1100100110100110", 30502 => "0110101110110110", 30503 => "1010110111001111", 30504 => "1111010110000110", 30505 => "0111010101110011", 30506 => "1001001000101001", 30507 => "1010010101100010", 30508 => "1001000110011101", 30509 => "0100111101100111", 30510 => "1000100010010101", 30511 => "1101111001010001", 30512 => "1000101010010010", 30513 => "1100000010111101", 30514 => "1000111101000010", 30515 => "1001011000001000", 30516 => "0010001100001110", 30517 => "1011110001110100", 30518 => "0110011110001110", 30519 => "0111101000110101", 30520 => "0010011010111110", 30521 => "1011110111111011", 30522 => "1011100011000011", 30523 => "0000010101001000", 30524 => "0011001001000001", 30525 => "1101011111100001", 30526 => "0101011110101000", 30527 => "1110000000001010", 30528 => "1001101010111100", 30529 => "1111110000001011", 30530 => "1101011101000111", 30531 => "0110011101001101", 30532 => "0101000001111010", 30533 => "0001100000101111", 30534 => "0011110001111010", 30535 => "1110001101111100", 30536 => "0000001010010111", 30537 => "0000110110111011", 30538 => "0011000001100000", 30539 => "1100001011101101", 30540 => "0000011111010110", 30541 => "0010001100000101", 30542 => "0010011000100110", 30543 => "1001111110011001", 30544 => "0000100010111110", 30545 => "1110111110010100", 30546 => "1111101110001011", 30547 => "0011010100011101", 30548 => "0010011000000101", 30549 => "0000011010101101", 30550 => "1000100110101000", 30551 => "1000110011111000", 30552 => "0100001011000111", 30553 => "0001100100111011", 30554 => "0000001101110000", 30555 => "1001010000101000", 30556 => "1111111101010001", 30557 => "0101010110001101", 30558 => "1111011000011000", 30559 => "0110000110011010", 30560 => "0110001110100100", 30561 => "0000000011001111", 30562 => "0101000000111000", 30563 => "0010110010111011", 30564 => "1011110011101110", 30565 => "1100010101110110", 30566 => "0010110000110100", 30567 => "1110001100011010", 30568 => "1101100001010001", 30569 => "1100001001110010", 30570 => "1110000011011110", 30571 => "0000110000100111", 30572 => "1101010001010000", 30573 => "0011111000100111", 30574 => "1101000000000011", 30575 => "0101111011100011", 30576 => "0000110000001100", 30577 => "0101011001011001", 30578 => "1110111110111101", 30579 => "0111010011100111", 30580 => "0001100111110011", 30581 => "0101000001100100", 30582 => "0111011001111011", 30583 => "1001001101111100", 30584 => "0000100001101110", 30585 => "1111101111110111", 30586 => "1011001001011001", 30587 => "1011011001011010", 30588 => "0101111001010100", 30589 => "0110001100011111", 30590 => "1000111000101101", 30591 => "1111110101011011", 30592 => "0000100100110111", 30593 => "1001010110110101", 30594 => "1010101101100110", 30595 => "1111111010011010", 30596 => "1110010100010011", 30597 => "1101100111010000", 30598 => "0001010000100101", 30599 => "0000110010011111", 30600 => "1010111010011010", 30601 => "1011001001110000", 30602 => "0001001101001101", 30603 => "1101110010011001", 30604 => "0101011110011000", 30605 => "1110011101101010", 30606 => "1110011001010000", 30607 => "1000010001110000", 30608 => "0010100000000011", 30609 => "0001110100110111", 30610 => "0111000000010010", 30611 => "1100111101011000", 30612 => "1000111000100011", 30613 => "0000001010100010", 30614 => "0000111011010111", 30615 => "1010110001110101", 30616 => "1011111010001100", 30617 => "1010001001100011", 30618 => "1100010010000000", 30619 => "1101110011001000", 30620 => "0100010001010000", 30621 => "1011000110111011", 30622 => "1000100101000100", 30623 => "0000100110110110", 30624 => "1011110101101110", 30625 => "1011100111101100", 30626 => "1111010010100110", 30627 => "1000001000001000", 30628 => "1110111001010010", 30629 => "0101010011011111", 30630 => "1001011010011110", 30631 => "1000001001001111", 30632 => "0010001111100001", 30633 => "1010100111110100", 30634 => "0101001011011000", 30635 => "0100100110010101", 30636 => "0001011011101111", 30637 => "1010110011100001", 30638 => "1010001101011101", 30639 => "0010010111111001", 30640 => "0000100101011011", 30641 => "1100110101010110", 30642 => "1101100010011110", 30643 => "1011111101011011", 30644 => "1111100011000100", 30645 => "0010010101111110", 30646 => "1010101000001001", 30647 => "0100000111111100", 30648 => "1111100111010111", 30649 => "1111101000001100", 30650 => "0100100010010111", 30651 => "1111000111000111", 30652 => "0101010111111000", 30653 => "1111001000010111", 30654 => "0100001011101100", 30655 => "1101111100000111", 30656 => "0110100101010011", 30657 => "1101111011101110", 30658 => "0001100000100101", 30659 => "1100000010101100", 30660 => "1110011110001110", 30661 => "1010000001110111", 30662 => "1110011110111111", 30663 => "0110001111011100", 30664 => "1101000100011110", 30665 => "0110010101001010", 30666 => "0010010111110000", 30667 => "1000001011001001", 30668 => "1000101000111010", 30669 => "0100110000110101", 30670 => "1101100110101001", 30671 => "0001001111001000", 30672 => "0101011110110010", 30673 => "0111111001100111", 30674 => "0110011101110101", 30675 => "1011101111111110", 30676 => "1000011001000010", 30677 => "0100100011000100", 30678 => "0101010100001100", 30679 => "0101010011101110", 30680 => "1111000101111000", 30681 => "1011100110010001", 30682 => "0011110101101010", 30683 => "0100110011010011", 30684 => "1010101101111101", 30685 => "1111100000000111", 30686 => "1010000110111110", 30687 => "1011011111011101", 30688 => "0101011100000101", 30689 => "1011011001000110", 30690 => "0101001001010011", 30691 => "1100110101000111", 30692 => "0110010101110110", 30693 => "0010011111010010", 30694 => "1100110001111011", 30695 => "1011000001011110", 30696 => "0110111011011110", 30697 => "0100111000000101", 30698 => "1100001001011001", 30699 => "0100001000000111", 30700 => "1101111001111000", 30701 => "0001101111011111", 30702 => "0011111001100010", 30703 => "0011111000101110", 30704 => "1011000001111110", 30705 => "0110111000000010", 30706 => "0110101011110010", 30707 => "0110001010111101", 30708 => "0101001001011111", 30709 => "1101100111001001", 30710 => "0000000110110110", 30711 => "0111010100100001", 30712 => "1111110100010001", 30713 => "1100101110111110", 30714 => "1100101001100110", 30715 => "0001011101111001", 30716 => "1100110111010100", 30717 => "1011100111111011", 30718 => "0110110111101101", 30719 => "1001100000000101", 30720 => "1111011010010111", 30721 => "1101011010000001", 30722 => "0010111111101100", 30723 => "0101111110010110", 30724 => "0100100011011100", 30725 => "0101000000000111", 30726 => "1101101101100101", 30727 => "1101101001100010", 30728 => "1000001100001001", 30729 => "0111101111101001", 30730 => "0100010010011010", 30731 => "1001111110001100", 30732 => "0110100001110000", 30733 => "1010100000101111", 30734 => "0101110011110000", 30735 => "0101011111000000", 30736 => "0001110111100011", 30737 => "0111110100010111", 30738 => "0010101101100001", 30739 => "1001011011001001", 30740 => "0110111111111001", 30741 => "1101111011011110", 30742 => "1100110001100010", 30743 => "0101010011010001", 30744 => "0110100110111110", 30745 => "1111111111100111", 30746 => "1100010111011101", 30747 => "0001011110101101", 30748 => "1001001110110110", 30749 => "1101101011001101", 30750 => "1100000101100001", 30751 => "1110110110011001", 30752 => "0111110010000110", 30753 => "0011010011001001", 30754 => "0110101010011101", 30755 => "0011100001110100", 30756 => "0000100111011000", 30757 => "0000110111011110", 30758 => "0101101010011001", 30759 => "1110001001000001", 30760 => "0101101110011101", 30761 => "1010100100100000", 30762 => "1011110000010011", 30763 => "0111010100111011", 30764 => "0101100001010110", 30765 => "0100010010111000", 30766 => "1000000001111111", 30767 => "1100001001010101", 30768 => "1101110101101100", 30769 => "1101111100100100", 30770 => "1101111001100011", 30771 => "1111011100110000", 30772 => "0011001011011011", 30773 => "0111101110010100", 30774 => "0100010011010110", 30775 => "0100111001011000", 30776 => "0101000110100000", 30777 => "0111000110011101", 30778 => "0101110011111010", 30779 => "1011101101101010", 30780 => "1010100111000100", 30781 => "0000110011010111", 30782 => "1101101100101101", 30783 => "1110011001010000", 30784 => "1111010011110101", 30785 => "1101001100100110", 30786 => "0111001100001001", 30787 => "0000111010000011", 30788 => "0110010101001001", 30789 => "0010101111001101", 30790 => "0011011110000110", 30791 => "0011000001110000", 30792 => "1110010101100101", 30793 => "0101101110011101", 30794 => "1100011001000101", 30795 => "1110101101110010", 30796 => "1001001110110011", 30797 => "1101100110010000", 30798 => "0011100100001001", 30799 => "1000010100111111", 30800 => "1101110100110111", 30801 => "0101100101110011", 30802 => "1111001100000101", 30803 => "1000101000010111", 30804 => "0001110101110100", 30805 => "1010101101110100", 30806 => "1000010100110101", 30807 => "0001110000111110", 30808 => "1100101101100100", 30809 => "1101000101110111", 30810 => "0101111111111010", 30811 => "1111010001010101", 30812 => "1101100110001011", 30813 => "0010101011001100", 30814 => "0001110010010110", 30815 => "0111001010010010", 30816 => "0001111100101001", 30817 => "0011111011110111", 30818 => "0101000111110101", 30819 => "0010110100100101", 30820 => "0011011101110010", 30821 => "1100100101110011", 30822 => "0010011010110000", 30823 => "0010000011010010", 30824 => "1011011010111111", 30825 => "0000001111110010", 30826 => "1110001000000001", 30827 => "1000110110001010", 30828 => "0001101000100000", 30829 => "1111101000111010", 30830 => "1010101011101110", 30831 => "0100101011111110", 30832 => "1011110100001010", 30833 => "1100001101110110", 30834 => "0100101110000101", 30835 => "1100110111011111", 30836 => "1010010011100101", 30837 => "0001000101010101", 30838 => "1101010001000000", 30839 => "0110010001001000", 30840 => "1101001110010111", 30841 => "1111101001011001", 30842 => "0110001111001000", 30843 => "0000001010111011", 30844 => "1000110011011111", 30845 => "1000100011001001", 30846 => "0010011100010100", 30847 => "0001000001000101", 30848 => "1111001001100110", 30849 => "0110111101111111", 30850 => "1100100001100101", 30851 => "1110111101001111", 30852 => "1001111011001100", 30853 => "1001111001001010", 30854 => "0011110100011110", 30855 => "1011110100110001", 30856 => "0000000010001100", 30857 => "0110011110111111", 30858 => "1000000010011010", 30859 => "1011001010001001", 30860 => "1011100101110110", 30861 => "1001010010001111", 30862 => "1111101100001001", 30863 => "0010011011100000", 30864 => "1100011101101101", 30865 => "1000110000010010", 30866 => "0100100110010111", 30867 => "0100100101001110", 30868 => "1110111011000111", 30869 => "0010000000111111", 30870 => "0110101110010100", 30871 => "0110110010011000", 30872 => "0110100110101100", 30873 => "0010000111010001", 30874 => "1010000011110101", 30875 => "0001000101110111", 30876 => "1111011010100010", 30877 => "1000111001111011", 30878 => "0011000101100011", 30879 => "0110011111111110", 30880 => "1001110011111000", 30881 => "1011011001010100", 30882 => "1110000111010001", 30883 => "0001111011001010", 30884 => "0001100001010100", 30885 => "1100101100110110", 30886 => "0000101111000010", 30887 => "0111000100001100", 30888 => "1010001101011010", 30889 => "1110010001111111", 30890 => "1100010001010000", 30891 => "0001110101000100", 30892 => "1111101101111100", 30893 => "0001101111001010", 30894 => "0011000110101110", 30895 => "0110000101101011", 30896 => "1110000101010111", 30897 => "0010111001101101", 30898 => "1111000110001101", 30899 => "0110010100000110", 30900 => "1100010011101100", 30901 => "0110100111010101", 30902 => "0110101100001111", 30903 => "0001101001001010", 30904 => "1110010000100110", 30905 => "0011111110000010", 30906 => "0100011011000000", 30907 => "0001110101010111", 30908 => "1100101011101101", 30909 => "0111110110011000", 30910 => "0101010010101110", 30911 => "1000010111010010", 30912 => "0000110100101100", 30913 => "1010110101000111", 30914 => "1010101111001010", 30915 => "1010111100111110", 30916 => "1101000011000001", 30917 => "0110001001111110", 30918 => "1001111000010011", 30919 => "1000100101100010", 30920 => "0001010111001010", 30921 => "1101111011100100", 30922 => "0111010111011001", 30923 => "0111100000100101", 30924 => "1001011001000000", 30925 => "1101100110100111", 30926 => "1000101000000010", 30927 => "1001101011001011", 30928 => "1001110101100111", 30929 => "0010011011101111", 30930 => "1110011111100110", 30931 => "0000000010110001", 30932 => "0010110010001111", 30933 => "0101101010110110", 30934 => "1001110001000100", 30935 => "1011010001010110", 30936 => "1110100111011101", 30937 => "1011010101111100", 30938 => "1110000010111101", 30939 => "1101110111111100", 30940 => "0100101010010001", 30941 => "1110100010011111", 30942 => "0101011000010111", 30943 => "1001111001111011", 30944 => "0110101101110110", 30945 => "1101000101101101", 30946 => "0001101001011111", 30947 => "1010101011101100", 30948 => "1110000010001011", 30949 => "0110010110101110", 30950 => "1010010101111100", 30951 => "1101110001000110", 30952 => "1000000111100110", 30953 => "0001110101110110", 30954 => "0101001011001111", 30955 => "0001011100010011", 30956 => "1011001000010100", 30957 => "1000010101001000", 30958 => "1001001010011011", 30959 => "1101101011001001", 30960 => "1011101100000010", 30961 => "0111000111111011", 30962 => "1000011100011100", 30963 => "1111011001100101", 30964 => "0111101111111111", 30965 => "1101100101111001", 30966 => "0110111000101011", 30967 => "1011001000101001", 30968 => "0010101111101100", 30969 => "1010010000101100", 30970 => "1110111001110010", 30971 => "0000101001111001", 30972 => "0110101010010100", 30973 => "0100011111000110", 30974 => "1100010111001111", 30975 => "0010111011111100", 30976 => "0100001010011101", 30977 => "1001101011110001", 30978 => "1011100001110000", 30979 => "1100001100000111", 30980 => "0100001011111000", 30981 => "0110000100110000", 30982 => "1110101111101001", 30983 => "1111001011001010", 30984 => "1010010100110000", 30985 => "1101010100101010", 30986 => "0101010111001110", 30987 => "0111000001100011", 30988 => "0111110000110010", 30989 => "0001011101010100", 30990 => "1100101100011001", 30991 => "1011100000111110", 30992 => "0001010101100011", 30993 => "0101001000011000", 30994 => "0011110100100101", 30995 => "0111011010101100", 30996 => "1110010101010000", 30997 => "0010001110101011", 30998 => "0111001001001010", 30999 => "1000100100000000", 31000 => "0100000100101101", 31001 => "1111101111100111", 31002 => "0111111001000101", 31003 => "1011010100110001", 31004 => "0011011010010000", 31005 => "1000000100000111", 31006 => "1010001101110011", 31007 => "0000011010000110", 31008 => "0100111101010001", 31009 => "0000111010101000", 31010 => "0011101001100010", 31011 => "0111001000011011", 31012 => "1100101111100100", 31013 => "1000011111110010", 31014 => "1011111000111101", 31015 => "0001110111010000", 31016 => "0111100111101101", 31017 => "0000011111110111", 31018 => "1111110101110110", 31019 => "1101001111000001", 31020 => "0010101000100111", 31021 => "0100010101010010", 31022 => "0000011101011110", 31023 => "1000101001111010", 31024 => "0110010101111110", 31025 => "0110101001100101", 31026 => "0110111010011000", 31027 => "1011100110011111", 31028 => "1011000101010110", 31029 => "0100101010000011", 31030 => "0010001111000111", 31031 => "0011111101100011", 31032 => "0101110101100011", 31033 => "0000111010011001", 31034 => "1001111010010010", 31035 => "1001010100100011", 31036 => "1100110100011001", 31037 => "1111101010111001", 31038 => "0101011000001001", 31039 => "1111101000011010", 31040 => "0001000100000001", 31041 => "0010001010110001", 31042 => "0111000000101100", 31043 => "1101000100100001", 31044 => "0000100101111000", 31045 => "1100001100101100", 31046 => "1010111001111100", 31047 => "0000001001001111", 31048 => "0110011001000001", 31049 => "0011011001001000", 31050 => "1110101001001001", 31051 => "0101101101000010", 31052 => "1110001100110111", 31053 => "0101101100011111", 31054 => "1110101110100010", 31055 => "1111111110011111", 31056 => "1110001110110111", 31057 => "1010011110100011", 31058 => "1000011010011010", 31059 => "0100001100111011", 31060 => "1111110101110011", 31061 => "0010000001011101", 31062 => "0011001001100110", 31063 => "0011011101000000", 31064 => "1101001110010010", 31065 => "1011101111101011", 31066 => "0100001011100000", 31067 => "1110010010010101", 31068 => "0000111010101101", 31069 => "1010111110110111", 31070 => "0000000101010100", 31071 => "0111101100110100", 31072 => "0011011111010001", 31073 => "1110111110011001", 31074 => "1111010001010111", 31075 => "0101011001001110", 31076 => "0110101000000010", 31077 => "0100110101010100", 31078 => "0101100010111100", 31079 => "1010100011000110", 31080 => "0110011000110010", 31081 => "0000011000001000", 31082 => "0001000010010000", 31083 => "1111000111100001", 31084 => "0010100110011111", 31085 => "1101111111110011", 31086 => "0100111100111000", 31087 => "1011010111101110", 31088 => "0100100101101110", 31089 => "0001000101010100", 31090 => "0010100100011110", 31091 => "1011110110100111", 31092 => "0101100000001010", 31093 => "0100100100101111", 31094 => "1111111001100011", 31095 => "1010110001001110", 31096 => "1100111111110111", 31097 => "0110111101011011", 31098 => "0100100010111010", 31099 => "1000010101001111", 31100 => "0100110111111100", 31101 => "0101011111101111", 31102 => "1011011111100111", 31103 => "1001000011000100", 31104 => "1101110011100100", 31105 => "0001101100000010", 31106 => "1001111010110001", 31107 => "0001010101101110", 31108 => "0111011000100100", 31109 => "0101001001110101", 31110 => "0111101100000011", 31111 => "0000000100011001", 31112 => "0111101001001000", 31113 => "0100011110000011", 31114 => "0111111000110011", 31115 => "1000101001101100", 31116 => "0010010100110110", 31117 => "0011100111101011", 31118 => "1001110111000011", 31119 => "0001111100001100", 31120 => "1001010010101000", 31121 => "0000001011011111", 31122 => "0001000010011110", 31123 => "0110001000011100", 31124 => "0011111011110010", 31125 => "0100011010011011", 31126 => "0100101000111111", 31127 => "1010111100000001", 31128 => "1001110011101000", 31129 => "1001011000001100", 31130 => "0101101000001010", 31131 => "1111110100010010", 31132 => "0001110100010010", 31133 => "1011001000000110", 31134 => "0001011110111100", 31135 => "0101001100001000", 31136 => "0010011100101100", 31137 => "0010011110101100", 31138 => "0010110011100110", 31139 => "0111010100010011", 31140 => "0101000001100001", 31141 => "0110010001101100", 31142 => "1010000000101001", 31143 => "1010000101010001", 31144 => "0111101110011001", 31145 => "1101001010000011", 31146 => "0001000101110011", 31147 => "0101011001111010", 31148 => "0101010011000100", 31149 => "1001100111101000", 31150 => "1110101100010100", 31151 => "0011001011001010", 31152 => "1101000101110011", 31153 => "1111100010101000", 31154 => "1111100010001010", 31155 => "0101110011011001", 31156 => "1101101111011010", 31157 => "1000010111111011", 31158 => "0000000100111000", 31159 => "0100001011010011", 31160 => "1110001010010011", 31161 => "1010110110110101", 31162 => "0111010010100001", 31163 => "0111011010010011", 31164 => "0011000001010000", 31165 => "0111110000000111", 31166 => "1110011010001001", 31167 => "1110110001101101", 31168 => "1110100001100011", 31169 => "1110100111000110", 31170 => "0111000110100100", 31171 => "1011000010100011", 31172 => "1000010001011110", 31173 => "0100101100100101", 31174 => "1111010001100001", 31175 => "1110011100100010", 31176 => "0110100101111101", 31177 => "1100011101100010", 31178 => "0000110010001110", 31179 => "1011010100101110", 31180 => "1000011011001011", 31181 => "1101011101100000", 31182 => "0010111010101000", 31183 => "1100101001100101", 31184 => "1010100010001111", 31185 => "1110010001100110", 31186 => "0010100100001100", 31187 => "1010110001010001", 31188 => "1110010110111010", 31189 => "0011100001001000", 31190 => "1111001000000110", 31191 => "0000000101111100", 31192 => "1101000111001010", 31193 => "1101100010000110", 31194 => "0110011101100001", 31195 => "1010110101111100", 31196 => "1001101010011110", 31197 => "0111110111001001", 31198 => "1100110011001000", 31199 => "1000001101111110", 31200 => "1011000101010001", 31201 => "0011100111011000", 31202 => "0001001101000111", 31203 => "1111100100101111", 31204 => "0000111001100010", 31205 => "0100011010111111", 31206 => "1110101101001000", 31207 => "1001111001100101", 31208 => "0101010010011100", 31209 => "1110110111011011", 31210 => "0011110111010101", 31211 => "1010111110100011", 31212 => "1101000111001011", 31213 => "1001101000011100", 31214 => "0100011010001101", 31215 => "0100001010101101", 31216 => "1001101100100110", 31217 => "1111000010000110", 31218 => "0100111001010011", 31219 => "1000000010010001", 31220 => "1010011000100010", 31221 => "0101011010000011", 31222 => "1011101100110101", 31223 => "0001010011100011", 31224 => "0100101010000010", 31225 => "0100100000111011", 31226 => "0011000100010101", 31227 => "1010111111101111", 31228 => "0100000001010000", 31229 => "0101000000010001", 31230 => "1101110111010111", 31231 => "1100000101100000", 31232 => "0111101101111110", 31233 => "1110011111010001", 31234 => "0111100010011111", 31235 => "1000011000010111", 31236 => "0111100111100001", 31237 => "0000101000101101", 31238 => "1010101001001011", 31239 => "1110010111111110", 31240 => "0010101011000111", 31241 => "0011101000101111", 31242 => "1111000100100001", 31243 => "1101010011101001", 31244 => "1100101011010100", 31245 => "0011010010011110", 31246 => "1010101100000000", 31247 => "0110000100000001", 31248 => "1101100100100000", 31249 => "1010010010100100", 31250 => "0010101010010111", 31251 => "1110110010101101", 31252 => "0100011001111101", 31253 => "0001001001010010", 31254 => "1101110111100100", 31255 => "1000001000110100", 31256 => "0011110110000101", 31257 => "1101111100110110", 31258 => "0111001011110100", 31259 => "1010000011000100", 31260 => "0010111111100101", 31261 => "1011100000101011", 31262 => "1101001001101101", 31263 => "1111000010100011", 31264 => "1100101101001011", 31265 => "0101100001111010", 31266 => "0011100010001001", 31267 => "1011010001011011", 31268 => "0010010001001111", 31269 => "1110011101001001", 31270 => "1100010110000110", 31271 => "0000000001110110", 31272 => "0111110111111101", 31273 => "0111010001000011", 31274 => "0001010011001000", 31275 => "1011001100001101", 31276 => "0001110010111100", 31277 => "1000101101001111", 31278 => "1101011011100100", 31279 => "0010000000000111", 31280 => "1111000100110111", 31281 => "1010000110110100", 31282 => "0110001110110110", 31283 => "1001111001110111", 31284 => "1101001010010001", 31285 => "1101100001110001", 31286 => "0010110011011010", 31287 => "0111110010111001", 31288 => "1100000110010111", 31289 => "1000100110101110", 31290 => "0000011100100001", 31291 => "1000011100111101", 31292 => "0000000001011000", 31293 => "0001110001111111", 31294 => "0110111101000001", 31295 => "1000110000000000", 31296 => "0000000001010000", 31297 => "1111101001010110", 31298 => "1000000010111111", 31299 => "0101001010111100", 31300 => "0001011011010100", 31301 => "0101110101001111", 31302 => "0000111010000011", 31303 => "1010011111001010", 31304 => "0000011110001001", 31305 => "1101111011000100", 31306 => "1001111111111110", 31307 => "0011100001100101", 31308 => "1111001000111110", 31309 => "0110111100001011", 31310 => "0111110110101100", 31311 => "1000010110010001", 31312 => "0110010000100110", 31313 => "1010011110000111", 31314 => "0110100111101000", 31315 => "0000001001010101", 31316 => "1111110101110000", 31317 => "0101011011010111", 31318 => "0111110100011111", 31319 => "1101011110111110", 31320 => "1101100111111111", 31321 => "1000100101101111", 31322 => "1101100011000101", 31323 => "1000111010100000", 31324 => "0100000001100000", 31325 => "0000011011101100", 31326 => "1111100100011001", 31327 => "0101000111111001", 31328 => "0100001101011010", 31329 => "0010000011110000", 31330 => "1100001100010011", 31331 => "1001110001001010", 31332 => "0011110101001010", 31333 => "1010000001000100", 31334 => "1101100000111100", 31335 => "1001011011100011", 31336 => "0100111011100011", 31337 => "0000100110001011", 31338 => "0011000000110011", 31339 => "0111000110010111", 31340 => "0110111000110101", 31341 => "0000111100000101", 31342 => "0010101011001100", 31343 => "1110001010001101", 31344 => "0000000100101000", 31345 => "1111011111011110", 31346 => "1111101001110000", 31347 => "0010000101000000", 31348 => "0100100110110011", 31349 => "1001111111000001", 31350 => "1001001001111100", 31351 => "1110101001101011", 31352 => "1111110000100100", 31353 => "1111100001010110", 31354 => "0101011001101001", 31355 => "0010001100101110", 31356 => "1000001101011101", 31357 => "0111110101111111", 31358 => "0100000110001011", 31359 => "1000111110000001", 31360 => "0111100101011011", 31361 => "1101001100000111", 31362 => "0101001100101000", 31363 => "0001011101001001", 31364 => "1110001111011110", 31365 => "0011011100110110", 31366 => "0111110111100101", 31367 => "1111000010011001", 31368 => "0011101001000100", 31369 => "0101010110010010", 31370 => "0101000101101110", 31371 => "0011011100001111", 31372 => "0010001111010111", 31373 => "0101100001001100", 31374 => "0010111010101110", 31375 => "1100010000000101", 31376 => "1110000100000010", 31377 => "1000000110010111", 31378 => "0110000010011100", 31379 => "0000001111110011", 31380 => "0100111011011111", 31381 => "0000000111111011", 31382 => "1011110110011011", 31383 => "0000001111011111", 31384 => "1111011001111100", 31385 => "0000001010000011", 31386 => "0010011011111000", 31387 => "1111110110110010", 31388 => "0000001101010000", 31389 => "1000000000110111", 31390 => "0100000010101101", 31391 => "1000011011100111", 31392 => "1101010101101101", 31393 => "0101101011010110", 31394 => "0001110010011100", 31395 => "1111101011000001", 31396 => "1001100101101001", 31397 => "0110001100011100", 31398 => "0000110110110010", 31399 => "0110101011000010", 31400 => "0001110000000111", 31401 => "1110100101111011", 31402 => "1011111011010010", 31403 => "0001101111011011", 31404 => "0011011000001011", 31405 => "0101101100000000", 31406 => "0100000010110000", 31407 => "0010100000001101", 31408 => "0001100100011111", 31409 => "0000100101011100", 31410 => "1011110010010010", 31411 => "0111101110110000", 31412 => "1001000110011001", 31413 => "0100010001011011", 31414 => "1000110000001011", 31415 => "1001001101101010", 31416 => "0110000001100101", 31417 => "1000101001001101", 31418 => "0000000101111001", 31419 => "0100110101000000", 31420 => "1001111001101101", 31421 => "0110001000001001", 31422 => "0100010111110101", 31423 => "0111101010110111", 31424 => "0010110011010110", 31425 => "1001110101010100", 31426 => "1111011001001100", 31427 => "1001010101100000", 31428 => "1000101111011100", 31429 => "0010111010101010", 31430 => "0110011001010000", 31431 => "1000001001110001", 31432 => "0000000001001000", 31433 => "1001101000010000", 31434 => "0110001101100100", 31435 => "1011001001101100", 31436 => "0001010100101111", 31437 => "1100101011111000", 31438 => "0001110001101100", 31439 => "0000111010100110", 31440 => "0111000001011000", 31441 => "0000001000001110", 31442 => "1111100010001110", 31443 => "0100000011011001", 31444 => "1110101001100011", 31445 => "1010011010001100", 31446 => "1001111111110111", 31447 => "0010011110000010", 31448 => "0010010101111000", 31449 => "0000101000100011", 31450 => "0010100011101001", 31451 => "1001100101101100", 31452 => "1111111110110111", 31453 => "1111100000010011", 31454 => "0001100111110101", 31455 => "0001010010011010", 31456 => "0001011100110100", 31457 => "0101101100010100", 31458 => "0110011100100010", 31459 => "0110101110100001", 31460 => "0101111001010010", 31461 => "0000011110011001", 31462 => "1010111010111111", 31463 => "0100111011011100", 31464 => "1011111110110011", 31465 => "1110101101111101", 31466 => "0000000111111011", 31467 => "1000011011011110", 31468 => "1101010001101100", 31469 => "0010101100101010", 31470 => "0000011110110111", 31471 => "1000110000100111", 31472 => "1010111111010110", 31473 => "0000111111110111", 31474 => "1001111110100101", 31475 => "0110110000001011", 31476 => "0110010101000010", 31477 => "0010100010010101", 31478 => "0010101011100000", 31479 => "1110010000000001", 31480 => "0100110100110101", 31481 => "0100101010001001", 31482 => "0001100111101100", 31483 => "0001101101000001", 31484 => "1011100010000111", 31485 => "1011001101010010", 31486 => "1100101000101101", 31487 => "1010001100110100", 31488 => "1110101101110101", 31489 => "0101000111011100", 31490 => "1010111111110011", 31491 => "0110110010000000", 31492 => "1100110010100011", 31493 => "1100101000101100", 31494 => "1100101001110101", 31495 => "0111010110111001", 31496 => "1001001101110101", 31497 => "0000110111010101", 31498 => "1000011101000001", 31499 => "0111010000101000", 31500 => "1110010000001000", 31501 => "0011111100000000", 31502 => "1100001000101110", 31503 => "0100100110101011", 31504 => "0000101100101010", 31505 => "1111111011101110", 31506 => "1000110010111011", 31507 => "1110100011010001", 31508 => "0110011000000011", 31509 => "1110010100011000", 31510 => "1110001101001110", 31511 => "1100001101100101", 31512 => "1100100100011101", 31513 => "0010110101100001", 31514 => "0111110101001101", 31515 => "0110100011001010", 31516 => "1101000111010111", 31517 => "0000100111110011", 31518 => "1110110110110101", 31519 => "1101000100111101", 31520 => "1101100111001100", 31521 => "1011011110110110", 31522 => "1110110011101000", 31523 => "0101110101100110", 31524 => "1101101010100010", 31525 => "0111101100100011", 31526 => "0011110111100000", 31527 => "0100100011001100", 31528 => "0100111010111001", 31529 => "1000110101011100", 31530 => "1110101000100100", 31531 => "0011101001100111", 31532 => "1111001100010010", 31533 => "0000100110110111", 31534 => "1110011101011111", 31535 => "1000000000101111", 31536 => "1010100000100111", 31537 => "1011101011000101", 31538 => "0110010111011011", 31539 => "1011001011110110", 31540 => "1001000110110100", 31541 => "0110000110011001", 31542 => "1001110000100100", 31543 => "1101111110110010", 31544 => "0110011001000001", 31545 => "0110011000000101", 31546 => "1011001000000000", 31547 => "0100101100010000", 31548 => "0000011011000000", 31549 => "1001000110010011", 31550 => "0010100100101100", 31551 => "0001001101001001", 31552 => "0001101100010101", 31553 => "0000000111100101", 31554 => "0100001100010101", 31555 => "1100101111000000", 31556 => "0110110001010101", 31557 => "1100101010011101", 31558 => "1001000001101011", 31559 => "0000000101011111", 31560 => "0111000110111110", 31561 => "0111100011010010", 31562 => "0010101001111000", 31563 => "0100110001111100", 31564 => "0100110011100011", 31565 => "0000011110110000", 31566 => "0110000010000001", 31567 => "1101000011100000", 31568 => "1000111001100110", 31569 => "1000011010010010", 31570 => "1101111000001011", 31571 => "1111100110111011", 31572 => "0110100011100110", 31573 => "0111010111011111", 31574 => "1111011011110101", 31575 => "1011000110000000", 31576 => "0011110100000101", 31577 => "1110100000011111", 31578 => "1111101001100110", 31579 => "1010110000001111", 31580 => "1001010111011101", 31581 => "1001000000110101", 31582 => "0101111110100100", 31583 => "0001100011101011", 31584 => "0100000011101111", 31585 => "0011010110110010", 31586 => "1011000000001111", 31587 => "1000110110011001", 31588 => "0000011001011111", 31589 => "0010010001000001", 31590 => "0011010110101111", 31591 => "1110111101011111", 31592 => "1011101110001001", 31593 => "1110010011110100", 31594 => "0011101011010011", 31595 => "0111110100010101", 31596 => "1010110011110100", 31597 => "1111011110100000", 31598 => "0101100000000011", 31599 => "0111000101010011", 31600 => "0110010010101101", 31601 => "0000000010110001", 31602 => "1110001010101110", 31603 => "0110011010001011", 31604 => "1100110011001101", 31605 => "0100100110110111", 31606 => "1110000001001010", 31607 => "0110001011010010", 31608 => "1100111110000001", 31609 => "0101101100110011", 31610 => "1110001000100101", 31611 => "1101000001010110", 31612 => "1101111010110101", 31613 => "1010101101111000", 31614 => "0000101110100100", 31615 => "1101110101110110", 31616 => "0010110011001111", 31617 => "0011000011001101", 31618 => "1001111001101101", 31619 => "0101100111101101", 31620 => "1101101010111000", 31621 => "1011010110011000", 31622 => "1000100110100001", 31623 => "1100111101001001", 31624 => "0111101101110101", 31625 => "0011101110100000", 31626 => "1100011111011111", 31627 => "0011000011101011", 31628 => "1100100111011010", 31629 => "1001101101010111", 31630 => "1100111101010000", 31631 => "1110110110111000", 31632 => "1000101001010011", 31633 => "0000101100111111", 31634 => "1101001100011101", 31635 => "1010001101111001", 31636 => "0110001001000010", 31637 => "1111001001011111", 31638 => "1001110000101110", 31639 => "0100111000001001", 31640 => "0010101001110111", 31641 => "0111001101101011", 31642 => "0010111110100111", 31643 => "0000011000000111", 31644 => "0110111001111111", 31645 => "0000100011100011", 31646 => "1001011100001000", 31647 => "0011011111100101", 31648 => "1111111010111110", 31649 => "1001101101100010", 31650 => "0110100111010001", 31651 => "1101101111111110", 31652 => "1100101101010100", 31653 => "0110111000001101", 31654 => "0001010001101110", 31655 => "0110011111001101", 31656 => "1100011001101100", 31657 => "1000101001010010", 31658 => "0011111110010111", 31659 => "0011100011000001", 31660 => "1110110010000111", 31661 => "1000110101110101", 31662 => "1000000100111001", 31663 => "1100101100001100", 31664 => "1001000011111010", 31665 => "1100100110110101", 31666 => "1011111001000101", 31667 => "1100000111001000", 31668 => "1010010000010000", 31669 => "1110011110001001", 31670 => "0001011110111110", 31671 => "1011110100110110", 31672 => "0110010100010011", 31673 => "1100110011011010", 31674 => "0100001011110000", 31675 => "0001001010110011", 31676 => "1011111100000110", 31677 => "0101100001001011", 31678 => "1011110111111110", 31679 => "1011011011000011", 31680 => "0011010001011011", 31681 => "1010011010110101", 31682 => "0010000110011110", 31683 => "0101010000000010", 31684 => "1111110010000011", 31685 => "1000011011011100", 31686 => "1000110011100101", 31687 => "1011000010100001", 31688 => "0101011111100001", 31689 => "1101100101101100", 31690 => "0110000001100001", 31691 => "0100101110011111", 31692 => "1111001011001011", 31693 => "1000110010000010", 31694 => "1100111110101000", 31695 => "0000111100001001", 31696 => "0100110110100110", 31697 => "0110100001111111", 31698 => "0001110100101111", 31699 => "1000101011010011", 31700 => "0001000011110010", 31701 => "0000101100110100", 31702 => "0111010101010000", 31703 => "0001001100010011", 31704 => "0001100011100001", 31705 => "0110001101011001", 31706 => "1010111111010110", 31707 => "0001111110100100", 31708 => "0000111000001100", 31709 => "0000011110100000", 31710 => "1101110000111000", 31711 => "1000111000101011", 31712 => "0001001001011110", 31713 => "0011101111010000", 31714 => "1110001011100011", 31715 => "0100100001000110", 31716 => "1111000010100100", 31717 => "0011010110000011", 31718 => "0100111111001110", 31719 => "1011010011110000", 31720 => "0101011001111010", 31721 => "1100100111101101", 31722 => "0000110001001110", 31723 => "1100000000011111", 31724 => "0000101110010100", 31725 => "1000001010001110", 31726 => "1100100110100011", 31727 => "1010010011100001", 31728 => "1111100101011110", 31729 => "0100100110011000", 31730 => "0100001010001001", 31731 => "0000111001101111", 31732 => "1101100011001001", 31733 => "0011110101110100", 31734 => "0010000100011000", 31735 => "0101110010101011", 31736 => "1101100001010100", 31737 => "0001001111110110", 31738 => "0010101001011101", 31739 => "1010001001000011", 31740 => "1100001110001001", 31741 => "1011001111001000", 31742 => "1011000010111010", 31743 => "0000000010001001", 31744 => "1011101001110111", 31745 => "0111110000110001", 31746 => "0111101000010001", 31747 => "1001010000111011", 31748 => "0001101000101111", 31749 => "0000110011000110", 31750 => "0110010100010100", 31751 => "0110001111001110", 31752 => "0001010100100100", 31753 => "0011111010101111", 31754 => "1111110011011011", 31755 => "1100111101000000", 31756 => "0101111011001110", 31757 => "1111010010110010", 31758 => "1011110101100101", 31759 => "1010001011101000", 31760 => "1110111111011011", 31761 => "1001010011001110", 31762 => "0111111000101101", 31763 => "0010100001001011", 31764 => "1100011001001011", 31765 => "0100010101100001", 31766 => "0111001011011010", 31767 => "1101000001111001", 31768 => "0000110111010011", 31769 => "0010110011011101", 31770 => "1010101101000111", 31771 => "1110011111110000", 31772 => "1010010001111101", 31773 => "0000110110000110", 31774 => "1101101011010110", 31775 => "0101011001111011", 31776 => "1001100100111111", 31777 => "0101011100101110", 31778 => "0011101100011101", 31779 => "1001110010111001", 31780 => "0100111110110100", 31781 => "0111101111011000", 31782 => "0001100000100100", 31783 => "1011011010001100", 31784 => "0010110100111011", 31785 => "1111111000111100", 31786 => "1111101101001010", 31787 => "0010001011010110", 31788 => "0111111011100000", 31789 => "0000110111101100", 31790 => "0111111000101101", 31791 => "1100011110001110", 31792 => "1101000001100010", 31793 => "0010100100001100", 31794 => "1111010010000010", 31795 => "1000101101010100", 31796 => "1011000110101100", 31797 => "0001010101100011", 31798 => "1011110011010101", 31799 => "0011100000010010", 31800 => "0100000011100011", 31801 => "0111001001100000", 31802 => "0010101111000101", 31803 => "0101101111111000", 31804 => "0001101011100001", 31805 => "0100110101101110", 31806 => "0100101100110111", 31807 => "1001000100000111", 31808 => "1100101001000000", 31809 => "0110100010101001", 31810 => "0010001100010111", 31811 => "1001100111001001", 31812 => "1011011110110011", 31813 => "1101100010111101", 31814 => "1111001010100010", 31815 => "0101011001101011", 31816 => "1100101011110000", 31817 => "0011111000101000", 31818 => "0101101110000101", 31819 => "0011000111000101", 31820 => "0011111111110110", 31821 => "0101111011101001", 31822 => "0100101100110100", 31823 => "0000110011110100", 31824 => "0101111001111110", 31825 => "0011110001101000", 31826 => "0010100001000110", 31827 => "1100110101010001", 31828 => "0100100111010000", 31829 => "0011111001110101", 31830 => "0010001100010001", 31831 => "0000110000110010", 31832 => "1010111000000000", 31833 => "0101110110110001", 31834 => "1111010011000010", 31835 => "1101010111110000", 31836 => "1001110101100101", 31837 => "0110000100011110", 31838 => "1000011100101000", 31839 => "1110011001011010", 31840 => "1111011100101001", 31841 => "0000001001001010", 31842 => "0011101101000000", 31843 => "0001011001001001", 31844 => "1101111010111001", 31845 => "1101110101100001", 31846 => "0111000100000011", 31847 => "1011111100001110", 31848 => "1011011000010011", 31849 => "1011100110100101", 31850 => "0100111101001110", 31851 => "1110101010011100", 31852 => "0111000110101101", 31853 => "1011001000010101", 31854 => "0111010101111101", 31855 => "1100000001000011", 31856 => "1111110011100011", 31857 => "0011000010111010", 31858 => "0100101011101001", 31859 => "0000111100001010", 31860 => "1110000110101000", 31861 => "1001001001110100", 31862 => "0000010101000011", 31863 => "1010000001101010", 31864 => "0010110010001000", 31865 => "1000001110100000", 31866 => "0100100101000000", 31867 => "0100101111100010", 31868 => "1001000001100010", 31869 => "1100001111101110", 31870 => "1011111001100011", 31871 => "0010101000001111", 31872 => "0101000100010011", 31873 => "1010111000100110", 31874 => "0100110111110101", 31875 => "1011110000101101", 31876 => "1010100111010011", 31877 => "1001101111011010", 31878 => "0000010001011011", 31879 => "0001111000011111", 31880 => "0101111101100000", 31881 => "1011101101111101", 31882 => "1110010101010110", 31883 => "1111101110000111", 31884 => "1111100101000000", 31885 => "0010101000110100", 31886 => "1101110000111011", 31887 => "0000100110011010", 31888 => "1010110111110010", 31889 => "0101111100111001", 31890 => "0100010100101110", 31891 => "1001011000100011", 31892 => "1011011001111011", 31893 => "1111001100011101", 31894 => "1100000011101010", 31895 => "0111010001010101", 31896 => "0001101110100011", 31897 => "1101111111010101", 31898 => "0011110010011010", 31899 => "0110010100111111", 31900 => "0011101001010111", 31901 => "0110010011100011", 31902 => "1110000110001011", 31903 => "0101101001101001", 31904 => "0010101100101100", 31905 => "1011010100000100", 31906 => "0010011010110001", 31907 => "0001000010111001", 31908 => "1101000011011100", 31909 => "1010000101111100", 31910 => "1110011001110011", 31911 => "0001001001100010", 31912 => "0101000011010110", 31913 => "0101100101111110", 31914 => "1010110111000001", 31915 => "1011111111110100", 31916 => "0111111010110101", 31917 => "1101100110100001", 31918 => "1011010011000000", 31919 => "1100110001100010", 31920 => "0110000110011101", 31921 => "0100101001001010", 31922 => "1000101010100011", 31923 => "1010100111001000", 31924 => "1010110111101101", 31925 => "1001001111101001", 31926 => "0000101001100100", 31927 => "1110000010011100", 31928 => "1110011000011001", 31929 => "1011100011011111", 31930 => "0001111011110101", 31931 => "1111111000001111", 31932 => "1111111000110000", 31933 => "0000011001101010", 31934 => "0000000001010001", 31935 => "1010100111101111", 31936 => "1111111101010111", 31937 => "1100010101111101", 31938 => "1111110010001111", 31939 => "0111110001010000", 31940 => "0111000011110101", 31941 => "1101110110110101", 31942 => "1001001111101001", 31943 => "1110000111100000", 31944 => "0001010011001111", 31945 => "0000110101101011", 31946 => "1010100000010101", 31947 => "0101011001000011", 31948 => "0001110000100011", 31949 => "1010001011000000", 31950 => "0001000110000011", 31951 => "1110111000111010", 31952 => "1100110010001111", 31953 => "1010101100111111", 31954 => "0110011001110011", 31955 => "1011000110011101", 31956 => "0101001110111010", 31957 => "0010011101101001", 31958 => "1111110011110110", 31959 => "0010011100101101", 31960 => "1000110100000101", 31961 => "1100010100000101", 31962 => "0000111011011110", 31963 => "0011101011100110", 31964 => "1000101010100101", 31965 => "1100101101000111", 31966 => "0011011011110000", 31967 => "1000110011110101", 31968 => "0010110001111010", 31969 => "0101110101011011", 31970 => "0100011100011001", 31971 => "0111100111101101", 31972 => "0110100000011100", 31973 => "1100011010101111", 31974 => "1111110010001111", 31975 => "1110100011111001", 31976 => "0010110010010110", 31977 => "1010101011011101", 31978 => "0011110110100110", 31979 => "1111010001010001", 31980 => "0011111000001010", 31981 => "0011001110010011", 31982 => "0001100001011011", 31983 => "0101110010000111", 31984 => "1011010010110000", 31985 => "1101101011110010", 31986 => "1000101100010000", 31987 => "1000001101111101", 31988 => "0111000100010101", 31989 => "1101010001011111", 31990 => "1111011110011101", 31991 => "0101000001010110", 31992 => "0100011111100110", 31993 => "0001010010010000", 31994 => "1011000101111000", 31995 => "1000100101010000", 31996 => "0100110011101000", 31997 => "1101010100001000", 31998 => "0011100010100110", 31999 => "0011111011000000", 32000 => "0011001000011010", 32001 => "0001000001001111", 32002 => "1111010010010101", 32003 => "1100100001101010", 32004 => "1111001101100011", 32005 => "0100101010111000", 32006 => "0100101001111101", 32007 => "1001011100100001", 32008 => "1000010111101010", 32009 => "0100101011011010", 32010 => "0010110001111011", 32011 => "0110001000101100", 32012 => "1110011100111101", 32013 => "1010000011011100", 32014 => "1110101000000011", 32015 => "1011101110111001", 32016 => "0010010110111100", 32017 => "0110100101000101", 32018 => "0110100110100100", 32019 => "1100001001111010", 32020 => "0000011100101111", 32021 => "0001100101011111", 32022 => "0010000001001100", 32023 => "0100000111011001", 32024 => "0100010101011111", 32025 => "0011001001000100", 32026 => "0111000101101100", 32027 => "1010011011110010", 32028 => "0010000010111010", 32029 => "1010000011000101", 32030 => "0101001010101010", 32031 => "1101110100010010", 32032 => "0111001011010100", 32033 => "0101100010111001", 32034 => "1111011110101101", 32035 => "0000111111110010", 32036 => "1011101001110000", 32037 => "1110101000101011", 32038 => "0110111100101100", 32039 => "1000100110110010", 32040 => "1111001110110000", 32041 => "0001111100011010", 32042 => "1000110111110101", 32043 => "0110111000111100", 32044 => "1010101001110000", 32045 => "1010000000010110", 32046 => "1010011100011011", 32047 => "1000111000101000", 32048 => "1001100100000001", 32049 => "0100101000000111", 32050 => "0110011100011101", 32051 => "0111000100011000", 32052 => "0010000101010001", 32053 => "0100000001010101", 32054 => "1100111001010101", 32055 => "0100110110101101", 32056 => "1110100111000110", 32057 => "1000010111101110", 32058 => "1010011000110111", 32059 => "1011001101110101", 32060 => "0010000111010111", 32061 => "1011110110011011", 32062 => "0101100000110001", 32063 => "0011101101010100", 32064 => "0010000010011011", 32065 => "1001011011111101", 32066 => "1011101111010000", 32067 => "1001010100010010", 32068 => "1001001111010110", 32069 => "1111000110101010", 32070 => "0001100101111111", 32071 => "1101011011100000", 32072 => "1011000111100111", 32073 => "1101010101111111", 32074 => "1011101100000111", 32075 => "0010100110011100", 32076 => "0100100000000011", 32077 => "1101000111011011", 32078 => "0001001011011101", 32079 => "1110100101100010", 32080 => "0101011010010001", 32081 => "0000010010111110", 32082 => "0101000101010110", 32083 => "0110110010110010", 32084 => "1100100010111000", 32085 => "1100111101111100", 32086 => "1011101100110000", 32087 => "1011101110111001", 32088 => "0100011000110101", 32089 => "0111111101110001", 32090 => "0000101010111000", 32091 => "0011001110110110", 32092 => "0100100111011100", 32093 => "0110010011000001", 32094 => "1110010000011111", 32095 => "1110101101100010", 32096 => "1010010111001000", 32097 => "0101000110100110", 32098 => "1111010010111000", 32099 => "1111110011010000", 32100 => "1011100001001100", 32101 => "1001001001101101", 32102 => "1010011101100101", 32103 => "0110111001010000", 32104 => "1000010111011010", 32105 => "0100100000111100", 32106 => "0100101100100011", 32107 => "0000101010101011", 32108 => "0011101101110010", 32109 => "0011001100000000", 32110 => "0100101101011010", 32111 => "1100100100111001", 32112 => "1000000110110001", 32113 => "0011000000010110", 32114 => "0000001011001001", 32115 => "0110000100010101", 32116 => "1110000111010101", 32117 => "0110101010001011", 32118 => "1001101011100100", 32119 => "1000010000100010", 32120 => "1000101001000011", 32121 => "0100000000110111", 32122 => "1010010010100001", 32123 => "1000011001010101", 32124 => "0001110100010010", 32125 => "1010010011000111", 32126 => "1011100100111100", 32127 => "1111001111000001", 32128 => "0011100010101111", 32129 => "0100111110100010", 32130 => "0010101011011010", 32131 => "0000010100110111", 32132 => "0011100101111111", 32133 => "0110011011000001", 32134 => "1110111111100111", 32135 => "1010111100101011", 32136 => "0100100010010011", 32137 => "0010001110110110", 32138 => "0110010000110011", 32139 => "0001010100001011", 32140 => "0001001110011011", 32141 => "0010111011101110", 32142 => "0001111001011110", 32143 => "1111010100101000", 32144 => "0111011111010101", 32145 => "0111011101011111", 32146 => "1010100011101111", 32147 => "0100110110000110", 32148 => "0011000011010101", 32149 => "1111011111001001", 32150 => "0000010011111000", 32151 => "1010011000001111", 32152 => "1101111000100010", 32153 => "0000000100101100", 32154 => "1001010101011000", 32155 => "1000100011111111", 32156 => "0011000110000001", 32157 => "1011011111011010", 32158 => "0101111000111101", 32159 => "1100001111111110", 32160 => "1001101001101100", 32161 => "0011111001010001", 32162 => "1101110100111110", 32163 => "0101000111010110", 32164 => "1010101010111010", 32165 => "1101100110100110", 32166 => "0111111111100100", 32167 => "0101000000011010", 32168 => "1110110011100111", 32169 => "1111101011111010", 32170 => "0001001010110000", 32171 => "1001011001000110", 32172 => "1000001001100011", 32173 => "1001011100111001", 32174 => "1011001010111011", 32175 => "1100111011101010", 32176 => "1011011101011110", 32177 => "1011111110100110", 32178 => "0100111100000110", 32179 => "1100100010110110", 32180 => "0101111000101100", 32181 => "0000010011100000", 32182 => "0011101100001110", 32183 => "1010000011110111", 32184 => "0110110110001010", 32185 => "1110100111011111", 32186 => "0110010000111010", 32187 => "0100101101100111", 32188 => "1101001100010110", 32189 => "0101001001011101", 32190 => "1111011010110010", 32191 => "0011010100111010", 32192 => "0000011100011110", 32193 => "0110010111100011", 32194 => "1001011110001010", 32195 => "1010011110100111", 32196 => "1001000000000011", 32197 => "1011011111100001", 32198 => "0011001111010010", 32199 => "0101111100001110", 32200 => "1101101001000101", 32201 => "0001010101111110", 32202 => "1110111000110010", 32203 => "0110000010111100", 32204 => "1111111111000000", 32205 => "0100010111011110", 32206 => "0001100001101001", 32207 => "1101100101100111", 32208 => "0101110011111011", 32209 => "1100010101011111", 32210 => "1100101001110100", 32211 => "1010001111000010", 32212 => "0001011000111010", 32213 => "1111110001011110", 32214 => "0101010110111011", 32215 => "0011110100101001", 32216 => "0001100010100010", 32217 => "0000100110101010", 32218 => "0100101011001111", 32219 => "1011111100011100", 32220 => "1011110110100000", 32221 => "1100000010111001", 32222 => "1100110100111100", 32223 => "1111101010010001", 32224 => "0000111010001111", 32225 => "1111110000001000", 32226 => "1101110011001010", 32227 => "0010100010111011", 32228 => "0011001011100001", 32229 => "1001000011001101", 32230 => "1110000001011000", 32231 => "0000001100000000", 32232 => "0001110001101001", 32233 => "1110100101100100", 32234 => "1111001010000111", 32235 => "0000011101001010", 32236 => "0101010111010100", 32237 => "0101000011100110", 32238 => "0111001101111100", 32239 => "0000101010010001", 32240 => "0011100001100010", 32241 => "1011000011000011", 32242 => "1110111101001101", 32243 => "1011011110100000", 32244 => "1110100110101111", 32245 => "1010001111000000", 32246 => "1101110010101101", 32247 => "0111110000001010", 32248 => "0011111000000100", 32249 => "0010000000001000", 32250 => "1110110010000111", 32251 => "1010001001111100", 32252 => "1101010011000000", 32253 => "0000100001010000", 32254 => "1110011001011000", 32255 => "1010000110111111", 32256 => "1010001010101111", 32257 => "0001101100011111", 32258 => "0010011100001000", 32259 => "0010110110011010", 32260 => "0001000000001111", 32261 => "1010111001100110", 32262 => "0100110100010010", 32263 => "0100011001001100", 32264 => "0100000101010111", 32265 => "0100010011001011", 32266 => "0100101011110100", 32267 => "0110010010001011", 32268 => "0010011111110110", 32269 => "0101000011100000", 32270 => "1110011011100000", 32271 => "1001000010000001", 32272 => "0010000110100010", 32273 => "0111100010000000", 32274 => "0100000100100011", 32275 => "0101111100101110", 32276 => "0101111000010111", 32277 => "1101101001110010", 32278 => "1111110110110101", 32279 => "0101101011010001", 32280 => "1110101111000001", 32281 => "0001000011111011", 32282 => "0101001100100111", 32283 => "1001000010110110", 32284 => "1000101010100101", 32285 => "1101101011100101", 32286 => "1010100111100110", 32287 => "1110010011000010", 32288 => "1010111101011011", 32289 => "1001101111010000", 32290 => "0100100100010110", 32291 => "1000001011101110", 32292 => "1010100010011111", 32293 => "1010000001101010", 32294 => "1000000100010111", 32295 => "1001010011001000", 32296 => "1100000010011110", 32297 => "1010100111000011", 32298 => "1111011011010101", 32299 => "0000000110100001", 32300 => "0111000001111110", 32301 => "1010100011000101", 32302 => "0001101110010100", 32303 => "1010100101111000", 32304 => "0001101111001000", 32305 => "0100111110110000", 32306 => "1111001111111000", 32307 => "1110011001101110", 32308 => "1000110100011101", 32309 => "0010100111111001", 32310 => "0100101111100011", 32311 => "1110010101011001", 32312 => "1111010010101110", 32313 => "1110110010110001", 32314 => "0010000100100101", 32315 => "0010000101101001", 32316 => "0011001111010001", 32317 => "0100011100100001", 32318 => "1011000110000100", 32319 => "0101110100100011", 32320 => "1011111101001011", 32321 => "0111001011000111", 32322 => "0000011101000011", 32323 => "0100110101100011", 32324 => "1110101111101001", 32325 => "1101000001100100", 32326 => "1011001110001010", 32327 => "0011010001110011", 32328 => "0010111011100011", 32329 => "0010010010101011", 32330 => "1011001100001010", 32331 => "1000000000010100", 32332 => "1000011111011010", 32333 => "1011000000101100", 32334 => "1100110101001100", 32335 => "1011001000101100", 32336 => "0111101011000000", 32337 => "1110110101011000", 32338 => "0010100100101000", 32339 => "0100101110100000", 32340 => "1001110001101011", 32341 => "0111001110010000", 32342 => "1011101101011100", 32343 => "1100001011111101", 32344 => "0100001101010010", 32345 => "1111001010100100", 32346 => "1011100101010000", 32347 => "1000101100010100", 32348 => "1100001011010110", 32349 => "0110111011100101", 32350 => "0000010011100001", 32351 => "0100000110100110", 32352 => "1100000001000011", 32353 => "0101100000110001", 32354 => "0011110100011101", 32355 => "1011010011000001", 32356 => "0111010101001001", 32357 => "1001111000010010", 32358 => "1101101010010010", 32359 => "1110111100110101", 32360 => "0101110001100111", 32361 => "0010010111101010", 32362 => "0101101000110110", 32363 => "1101010000010010", 32364 => "0000101111100000", 32365 => "1011110000110011", 32366 => "1000101101111101", 32367 => "0111011001000011", 32368 => "0111100010110010", 32369 => "1001101001111011", 32370 => "0011001011010100", 32371 => "0000110001101101", 32372 => "0011111010110010", 32373 => "1010010101000110", 32374 => "1000010100111111", 32375 => "1001111101111101", 32376 => "1110011001100111", 32377 => "0011100010010011", 32378 => "1001111101111101", 32379 => "1011100011100110", 32380 => "1011110101010011", 32381 => "1011011110110100", 32382 => "0011010010001101", 32383 => "0001001011110010", 32384 => "0100000000100001", 32385 => "1100100000011101", 32386 => "0011001100111110", 32387 => "1101010001001010", 32388 => "1011100010000000", 32389 => "1100010010010101", 32390 => "1111000101110111", 32391 => "1110101101111100", 32392 => "1110101111110111", 32393 => "0100000101011100", 32394 => "1001111111000110", 32395 => "0010101100010101", 32396 => "1100110111100100", 32397 => "1010101000000111", 32398 => "1101100111101101", 32399 => "1101000001011111", 32400 => "0001011011001101", 32401 => "1000100000010101", 32402 => "0100001000000010", 32403 => "1111110100101000", 32404 => "1001001111111000", 32405 => "1010111000100011", 32406 => "1101111100001101", 32407 => "0011101001011101", 32408 => "0100101010010101", 32409 => "0010111011111110", 32410 => "1000111101000110", 32411 => "1101111010010111", 32412 => "0001011101011100", 32413 => "1101010101010111", 32414 => "1101101001000001", 32415 => "1100110001010010", 32416 => "1011110111111111", 32417 => "0101000000011011", 32418 => "1000100001101111", 32419 => "1110000010101000", 32420 => "0001101001000101", 32421 => "0011010110010110", 32422 => "0100000000000000", 32423 => "0110100011100100", 32424 => "0010010100100110", 32425 => "1100100001101011", 32426 => "1101001010100010", 32427 => "0110001000001100", 32428 => "0100010111001001", 32429 => "0000101101010001", 32430 => "0000011000001011", 32431 => "1111010101001100", 32432 => "1000010111000010", 32433 => "0011111101011100", 32434 => "1110101111001110", 32435 => "0101011001110101", 32436 => "1000010010100110", 32437 => "1010011111100010", 32438 => "1101001001000001", 32439 => "1001010111101001", 32440 => "0111000000110011", 32441 => "0011101100000010", 32442 => "0101100100100100", 32443 => "0100000000010101", 32444 => "0110100001011100", 32445 => "1111001011011101", 32446 => "1110000000010001", 32447 => "1001100100011001", 32448 => "1110011010001111", 32449 => "0001100010111000", 32450 => "0111101001010001", 32451 => "0000111011100010", 32452 => "0000011010001110", 32453 => "0110100011000010", 32454 => "0011011011001000", 32455 => "0111010000101001", 32456 => "0101001100000001", 32457 => "0000011001110100", 32458 => "1000010011100010", 32459 => "0011100100111001", 32460 => "0101001101001101", 32461 => "1011101001000011", 32462 => "1001011010100010", 32463 => "0011110000001010", 32464 => "0111101111011110", 32465 => "1111001010111010", 32466 => "1001100110111010", 32467 => "1110101110100010", 32468 => "0010110100001011", 32469 => "1111110101011010", 32470 => "0101000101101001", 32471 => "0111011000110100", 32472 => "0000010101110000", 32473 => "0110100010011101", 32474 => "1100110101011110", 32475 => "0100011000000101", 32476 => "0010010001110000", 32477 => "1101000100110101", 32478 => "1110100010101010", 32479 => "1100011010010010", 32480 => "1111000110110110", 32481 => "1110010100001111", 32482 => "0110110010100001", 32483 => "1110101001100000", 32484 => "1010000100000000", 32485 => "1011001100100111", 32486 => "1001101010010001", 32487 => "1111000011101110", 32488 => "1000011010100101", 32489 => "0110000111001101", 32490 => "0101111010001001", 32491 => "0001101000000000", 32492 => "1101110101110110", 32493 => "0110101000100100", 32494 => "1010101011011001", 32495 => "0010011110001001", 32496 => "1100100000010100", 32497 => "1011000101111011", 32498 => "1110011000110011", 32499 => "0000011111001011", 32500 => "1011110101110011", 32501 => "0110010101011110", 32502 => "1011000100001000", 32503 => "0101000111100110", 32504 => "1011101101100001", 32505 => "1100010111000100", 32506 => "0010011000011010", 32507 => "1001010010100001", 32508 => "0010000010110011", 32509 => "0000110000110111", 32510 => "0100011001011001", 32511 => "1100010000010010", 32512 => "1111110011110010", 32513 => "0110010101110011", 32514 => "0111011001011101", 32515 => "1101011011011001", 32516 => "1011101101101011", 32517 => "0100010010110011", 32518 => "0100101111110010", 32519 => "1001001110011001", 32520 => "0111000101001111", 32521 => "0000001101110110", 32522 => "0101000010110110", 32523 => "0001000111111101", 32524 => "0011101111010101", 32525 => "0000111111100110", 32526 => "1110000100111000", 32527 => "1010100001011011", 32528 => "0010001100000010", 32529 => "0100010010100110", 32530 => "1101011000100000", 32531 => "0011011011001001", 32532 => "0000000011111101", 32533 => "0011101101101111", 32534 => "1010110001011010", 32535 => "0101110101010100", 32536 => "0010100100011011", 32537 => "0010010011100010", 32538 => "1001111001111110", 32539 => "1010111001010000", 32540 => "1101100101011000", 32541 => "0011001111110110", 32542 => "0000110101101100", 32543 => "0101011110001010", 32544 => "0111100101000100", 32545 => "0001101011001010", 32546 => "1100011000100100", 32547 => "0001011001101111", 32548 => "1101001010100101", 32549 => "0011010101011111", 32550 => "0000110010100000", 32551 => "1001110110011011", 32552 => "0100101111010110", 32553 => "1101101101101111", 32554 => "1010110011101111", 32555 => "0111100011110001", 32556 => "1001100101000111", 32557 => "0000101010011110", 32558 => "0000110111010011", 32559 => "1011101101010101", 32560 => "1101001000111010", 32561 => "1001111001000000", 32562 => "0011001111110100", 32563 => "0110100010000110", 32564 => "1000101110110110", 32565 => "0010001011110100", 32566 => "1010100010100000", 32567 => "0111101100011111", 32568 => "0000010000111011", 32569 => "1001111001101100", 32570 => "1001101101101001", 32571 => "1010011011000100", 32572 => "1110101110100011", 32573 => "1011000111011000", 32574 => "1110110001010100", 32575 => "1110111111001001", 32576 => "0001110001101111", 32577 => "1010000101111011", 32578 => "1110001000100010", 32579 => "1011100110100110", 32580 => "0111010001011111", 32581 => "1001010001100010", 32582 => "0001100111101011", 32583 => "0111110111011010", 32584 => "0111000100110111", 32585 => "0011100101101000", 32586 => "1111110001011111", 32587 => "0110110000010101", 32588 => "1100010101010111", 32589 => "0010001110011000", 32590 => "0100101010001111", 32591 => "1111010000110010", 32592 => "1010011010010011", 32593 => "0011011000011100", 32594 => "1001001111110010", 32595 => "0110110111101101", 32596 => "0000100111010100", 32597 => "1100101110101111", 32598 => "0010001111101110", 32599 => "1110110010011110", 32600 => "1000100000110100", 32601 => "1110110000001101", 32602 => "1001011011001000", 32603 => "1001110100110011", 32604 => "1111000011100010", 32605 => "0001100000010010", 32606 => "0000011110011100", 32607 => "0101111100101011", 32608 => "1100000010100101", 32609 => "0101011000010100", 32610 => "1110101010110110", 32611 => "1101011010110110", 32612 => "1101000011110000", 32613 => "0101010110100000", 32614 => "0110000101100001", 32615 => "0100100010000100", 32616 => "0111101100010101", 32617 => "1010110100110011", 32618 => "0100001110111011", 32619 => "1101101111011111", 32620 => "0011001110011111", 32621 => "0010110110100011", 32622 => "1000010101010001", 32623 => "1101111001010010", 32624 => "1011001011000101", 32625 => "0111101011111111", 32626 => "0010011101110001", 32627 => "0000011000111011", 32628 => "1111000100010111", 32629 => "1111000110111000", 32630 => "0010110010100100", 32631 => "1010010110001010", 32632 => "0000000111010011", 32633 => "1110001000001011", 32634 => "0100001000010001", 32635 => "1001101100100000", 32636 => "1010011111011001", 32637 => "0110001000010001", 32638 => "1001011011011011", 32639 => "1011101000100000", 32640 => "0001000110001011", 32641 => "1101111011001101", 32642 => "1011010101001111", 32643 => "1010111101000111", 32644 => "1101011101001010", 32645 => "1000101010100101", 32646 => "1111111010110001", 32647 => "0101101110000001", 32648 => "0001011111011001", 32649 => "1100111011110001", 32650 => "1000111010111001", 32651 => "0101000101101101", 32652 => "1011111000101110", 32653 => "0101110010100010", 32654 => "1110010001100110", 32655 => "1110111111011000", 32656 => "1101100011111001", 32657 => "1111000110101100", 32658 => "0010110101000010", 32659 => "0011111110000100", 32660 => "0110100010000010", 32661 => "1011010101000110", 32662 => "0100100110011110", 32663 => "1001000011111000", 32664 => "1111101111101100", 32665 => "0110011100100110", 32666 => "0010111000001110", 32667 => "0111100100010100", 32668 => "0101100111011011", 32669 => "0000000010111110", 32670 => "0110000001010101", 32671 => "0010000000000111", 32672 => "0000001001110000", 32673 => "1100000001111011", 32674 => "0110001101100010", 32675 => "0001100101010010", 32676 => "0011011100101111", 32677 => "0100111110100000", 32678 => "0101000111100010", 32679 => "1111111000010000", 32680 => "0110110000100111", 32681 => "1010111011110001", 32682 => "0000011011100001", 32683 => "1110011100110101", 32684 => "0010100101111110", 32685 => "0111011011100101", 32686 => "1001110001100101", 32687 => "0000010110100001", 32688 => "1101100110110101", 32689 => "0101110010010101", 32690 => "0100110001001011", 32691 => "0001010010110001", 32692 => "0101001100100110", 32693 => "0010011110001111", 32694 => "1011010100010010", 32695 => "0101110110111011", 32696 => "1010001101000111", 32697 => "0010011111111000", 32698 => "1010100110000101", 32699 => "0100000111100101", 32700 => "1110100011001101", 32701 => "0010111001100110", 32702 => "1001001101100000", 32703 => "0110111100010110", 32704 => "1011111101010000", 32705 => "1010000010000000", 32706 => "1101110001001100", 32707 => "0001000010110100", 32708 => "1101111011111111", 32709 => "1110100010000101", 32710 => "0101010101010110", 32711 => "1101111101110111", 32712 => "1100100010010110", 32713 => "1001111101100110", 32714 => "1100000011010011", 32715 => "1110111110110101", 32716 => "0000101010011010", 32717 => "1001000101100111", 32718 => "1010111110000100", 32719 => "1110111100010110", 32720 => "1011000111100101", 32721 => "0100111010001000", 32722 => "0101111000111110", 32723 => "0010101101010101", 32724 => "1010101010111110", 32725 => "1100011011111111", 32726 => "1011111100000001", 32727 => "0001000000011100", 32728 => "1100100111111001", 32729 => "1101000010001110", 32730 => "1000010000000100", 32731 => "0101111001100011", 32732 => "0110101100101100", 32733 => "1001101001110101", 32734 => "1100101101001100", 32735 => "1100001011110110", 32736 => "1010001100100101", 32737 => "0001101010101111", 32738 => "1010101001011001", 32739 => "0110100001110000", 32740 => "0110100111100111", 32741 => "1110111001010111", 32742 => "0011100101100011", 32743 => "0101011011010100", 32744 => "1000110000011110", 32745 => "1001101001000100", 32746 => "0001010110100100", 32747 => "1101000111110010", 32748 => "1010000111000000", 32749 => "1010111110011010", 32750 => "0011010000001110", 32751 => "0010110000000110", 32752 => "1100000010110101", 32753 => "0010100010101111", 32754 => "0000101001110000", 32755 => "0000100010110011", 32756 => "0111001010101011", 32757 => "1010111010110100", 32758 => "1010000111011110", 32759 => "0001101100001100", 32760 => "1110001001011010", 32761 => "0110001001001001", 32762 => "0001010010011101", 32763 => "0111011101011100", 32764 => "1001101010100011", 32765 => "0001110111010011", 32766 => "1010111011001111", 32767 => "1000100100011000");
BEGIN
  data_out <= ROM(to_integer(unsigned(address)));
END ARCHITECTURE;
