LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY rom IS
  PORT (
    address : IN STD_ULOGIC_VECTOR(14 DOWNTO 0);
    data_out : OUT STD_ULOGIC_VECTOR(15 DOWNTO 0));
END ENTITY;

ARCHITECTURE behavioural OF rom IS
  TYPE ROM_type IS ARRAY (0 TO 32767) OF STD_ULOGIC_VECTOR(15 DOWNTO 0);
  CONSTANT ROM : ROM_type := (0 => "0100000000000000", 1 => "1110101010001000", 2 => "0000000000000010", 3 => "1110101010001000", 4 => "0000000000000001", 5 => "1110101010001000", 6 => "0000000000000000", 7 => "1110101010001000", 8 => "0000000000000000", 9 => "1111110111001000", 10 => "0000000001100011", 11 => "1110110000010000", 12 => "0000000000000110", 13 => "1111000111000100", 14 => "0000000000000001", 15 => "1111110111001000", 16 => "0000001111101000", 17 => "1110110000010000", 18 => "0000000000000100", 19 => "1111000111000100", 20 => "0000000000000010", 21 => "1111110111001000", 22 => "0000001111101000", 23 => "1110110000010000", 24 => "0000000000000010", 25 => "1111000111000100", 26 => "0100000000000000", 27 => "1110111111001000", 28 => "0000000000000010", 29 => "1110101010001000", 30 => "0000000000000001", 31 => "1110101010001000", 32 => "0000000000000000", 33 => "1110101010001000", 34 => "0000000000000000", 35 => "1111110111001000", 36 => "0000000001100011", 37 => "1110110000010000", 38 => "0000000000100000", 39 => "1111000111000100", 40 => "0000000000000001", 41 => "1111110111001000", 42 => "0000001111101000", 43 => "1110110000010000", 44 => "0000000000011110", 45 => "1111000111000100", 46 => "0000000000000010", 47 => "1111110111001000", 48 => "0000001111101000", 49 => "1110110000010000", 50 => "0000000000011100", 51 => "1111000111000100", 52 => "0000000000000000", 53 => "1110101010000111", 54 => "0000000000000000", 55 => "0000000000000000", 56 => "0000000000000000", 57 => "0000000000000000", 58 => "0000000000000000", 59 => "0000000000000000", 60 => "0000000000000000", 61 => "0000000000000000", 62 => "0000000000000000", 63 => "0000000000000000", 64 => "0000000000000000", 65 => "0000000000000000", 66 => "0000000000000000", 67 => "0000000000000000", 68 => "0000000000000000", 69 => "0000000000000000", 70 => "0000000000000000", 71 => "0000000000000000", 72 => "0000000000000000", 73 => "0000000000000000", 74 => "0000000000000000", 75 => "0000000000000000", 76 => "0000000000000000", 77 => "0000000000000000", 78 => "0000000000000000", 79 => "0000000000000000", 80 => "0000000000000000", 81 => "0000000000000000", 82 => "0000000000000000", 83 => "0000000000000000", 84 => "0000000000000000", 85 => "0000000000000000", 86 => "0000000000000000", 87 => "0000000000000000", 88 => "0000000000000000", 89 => "0000000000000000", 90 => "0000000000000000", 91 => "0000000000000000", 92 => "0000000000000000", 93 => "0000000000000000", 94 => "0000000000000000", 95 => "0000000000000000", 96 => "0000000000000000", 97 => "0000000000000000", 98 => "0000000000000000", 99 => "0000000000000000", 100 => "0000000000000000", 101 => "0000000000000000", 102 => "0000000000000000", 103 => "0000000000000000", 104 => "0000000000000000", 105 => "0000000000000000", 106 => "0000000000000000", 107 => "0000000000000000", 108 => "0000000000000000", 109 => "0000000000000000", 110 => "0000000000000000", 111 => "0000000000000000", 112 => "0000000000000000", 113 => "0000000000000000", 114 => "0000000000000000", 115 => "0000000000000000", 116 => "0000000000000000", 117 => "0000000000000000", 118 => "0000000000000000", 119 => "0000000000000000", 120 => "0000000000000000", 121 => "0000000000000000", 122 => "0000000000000000", 123 => "0000000000000000", 124 => "0000000000000000", 125 => "0000000000000000", 126 => "0000000000000000", 127 => "0000000000000000", 128 => "0000000000000000", 129 => "0000000000000000", 130 => "0000000000000000", 131 => "0000000000000000", 132 => "0000000000000000", 133 => "0000000000000000", 134 => "0000000000000000", 135 => "0000000000000000", 136 => "0000000000000000", 137 => "0000000000000000", 138 => "0000000000000000", 139 => "0000000000000000", 140 => "0000000000000000", 141 => "0000000000000000", 142 => "0000000000000000", 143 => "0000000000000000", 144 => "0000000000000000", 145 => "0000000000000000", 146 => "0000000000000000", 147 => "0000000000000000", 148 => "0000000000000000", 149 => "0000000000000000", 150 => "0000000000000000", 151 => "0000000000000000", 152 => "0000000000000000", 153 => "0000000000000000", 154 => "0000000000000000", 155 => "0000000000000000", 156 => "0000000000000000", 157 => "0000000000000000", 158 => "0000000000000000", 159 => "0000000000000000", 160 => "0000000000000000", 161 => "0000000000000000", 162 => "0000000000000000", 163 => "0000000000000000", 164 => "0000000000000000", 165 => "0000000000000000", 166 => "0000000000000000", 167 => "0000000000000000", 168 => "0000000000000000", 169 => "0000000000000000", 170 => "0000000000000000", 171 => "0000000000000000", 172 => "0000000000000000", 173 => "0000000000000000", 174 => "0000000000000000", 175 => "0000000000000000", 176 => "0000000000000000", 177 => "0000000000000000", 178 => "0000000000000000", 179 => "0000000000000000", 180 => "0000000000000000", 181 => "0000000000000000", 182 => "0000000000000000", 183 => "0000000000000000", 184 => "0000000000000000", 185 => "0000000000000000", 186 => "0000000000000000", 187 => "0000000000000000", 188 => "0000000000000000", 189 => "0000000000000000", 190 => "0000000000000000", 191 => "0000000000000000", 192 => "0000000000000000", 193 => "0000000000000000", 194 => "0000000000000000", 195 => "0000000000000000", 196 => "0000000000000000", 197 => "0000000000000000", 198 => "0000000000000000", 199 => "0000000000000000", 200 => "0000000000000000", 201 => "0000000000000000", 202 => "0000000000000000", 203 => "0000000000000000", 204 => "0000000000000000", 205 => "0000000000000000", 206 => "0000000000000000", 207 => "0000000000000000", 208 => "0000000000000000", 209 => "0000000000000000", 210 => "0000000000000000", 211 => "0000000000000000", 212 => "0000000000000000", 213 => "0000000000000000", 214 => "0000000000000000", 215 => "0000000000000000", 216 => "0000000000000000", 217 => "0000000000000000", 218 => "0000000000000000", 219 => "0000000000000000", 220 => "0000000000000000", 221 => "0000000000000000", 222 => "0000000000000000", 223 => "0000000000000000", 224 => "0000000000000000", 225 => "0000000000000000", 226 => "0000000000000000", 227 => "0000000000000000", 228 => "0000000000000000", 229 => "0000000000000000", 230 => "0000000000000000", 231 => "0000000000000000", 232 => "0000000000000000", 233 => "0000000000000000", 234 => "0000000000000000", 235 => "0000000000000000", 236 => "0000000000000000", 237 => "0000000000000000", 238 => "0000000000000000", 239 => "0000000000000000", 240 => "0000000000000000", 241 => "0000000000000000", 242 => "0000000000000000", 243 => "0000000000000000", 244 => "0000000000000000", 245 => "0000000000000000", 246 => "0000000000000000", 247 => "0000000000000000", 248 => "0000000000000000", 249 => "0000000000000000", 250 => "0000000000000000", 251 => "0000000000000000", 252 => "0000000000000000", 253 => "0000000000000000", 254 => "0000000000000000", 255 => "0000000000000000", 256 => "0000000000000000", 257 => "0000000000000000", 258 => "0000000000000000", 259 => "0000000000000000", 260 => "0000000000000000", 261 => "0000000000000000", 262 => "0000000000000000", 263 => "0000000000000000", 264 => "0000000000000000", 265 => "0000000000000000", 266 => "0000000000000000", 267 => "0000000000000000", 268 => "0000000000000000", 269 => "0000000000000000", 270 => "0000000000000000", 271 => "0000000000000000", 272 => "0000000000000000", 273 => "0000000000000000", 274 => "0000000000000000", 275 => "0000000000000000", 276 => "0000000000000000", 277 => "0000000000000000", 278 => "0000000000000000", 279 => "0000000000000000", 280 => "0000000000000000", 281 => "0000000000000000", 282 => "0000000000000000", 283 => "0000000000000000", 284 => "0000000000000000", 285 => "0000000000000000", 286 => "0000000000000000", 287 => "0000000000000000", 288 => "0000000000000000", 289 => "0000000000000000", 290 => "0000000000000000", 291 => "0000000000000000", 292 => "0000000000000000", 293 => "0000000000000000", 294 => "0000000000000000", 295 => "0000000000000000", 296 => "0000000000000000", 297 => "0000000000000000", 298 => "0000000000000000", 299 => "0000000000000000", 300 => "0000000000000000", 301 => "0000000000000000", 302 => "0000000000000000", 303 => "0000000000000000", 304 => "0000000000000000", 305 => "0000000000000000", 306 => "0000000000000000", 307 => "0000000000000000", 308 => "0000000000000000", 309 => "0000000000000000", 310 => "0000000000000000", 311 => "0000000000000000", 312 => "0000000000000000", 313 => "0000000000000000", 314 => "0000000000000000", 315 => "0000000000000000", 316 => "0000000000000000", 317 => "0000000000000000", 318 => "0000000000000000", 319 => "0000000000000000", 320 => "0000000000000000", 321 => "0000000000000000", 322 => "0000000000000000", 323 => "0000000000000000", 324 => "0000000000000000", 325 => "0000000000000000", 326 => "0000000000000000", 327 => "0000000000000000", 328 => "0000000000000000", 329 => "0000000000000000", 330 => "0000000000000000", 331 => "0000000000000000", 332 => "0000000000000000", 333 => "0000000000000000", 334 => "0000000000000000", 335 => "0000000000000000", 336 => "0000000000000000", 337 => "0000000000000000", 338 => "0000000000000000", 339 => "0000000000000000", 340 => "0000000000000000", 341 => "0000000000000000", 342 => "0000000000000000", 343 => "0000000000000000", 344 => "0000000000000000", 345 => "0000000000000000", 346 => "0000000000000000", 347 => "0000000000000000", 348 => "0000000000000000", 349 => "0000000000000000", 350 => "0000000000000000", 351 => "0000000000000000", 352 => "0000000000000000", 353 => "0000000000000000", 354 => "0000000000000000", 355 => "0000000000000000", 356 => "0000000000000000", 357 => "0000000000000000", 358 => "0000000000000000", 359 => "0000000000000000", 360 => "0000000000000000", 361 => "0000000000000000", 362 => "0000000000000000", 363 => "0000000000000000", 364 => "0000000000000000", 365 => "0000000000000000", 366 => "0000000000000000", 367 => "0000000000000000", 368 => "0000000000000000", 369 => "0000000000000000", 370 => "0000000000000000", 371 => "0000000000000000", 372 => "0000000000000000", 373 => "0000000000000000", 374 => "0000000000000000", 375 => "0000000000000000", 376 => "0000000000000000", 377 => "0000000000000000", 378 => "0000000000000000", 379 => "0000000000000000", 380 => "0000000000000000", 381 => "0000000000000000", 382 => "0000000000000000", 383 => "0000000000000000", 384 => "0000000000000000", 385 => "0000000000000000", 386 => "0000000000000000", 387 => "0000000000000000", 388 => "0000000000000000", 389 => "0000000000000000", 390 => "0000000000000000", 391 => "0000000000000000", 392 => "0000000000000000", 393 => "0000000000000000", 394 => "0000000000000000", 395 => "0000000000000000", 396 => "0000000000000000", 397 => "0000000000000000", 398 => "0000000000000000", 399 => "0000000000000000", 400 => "0000000000000000", 401 => "0000000000000000", 402 => "0000000000000000", 403 => "0000000000000000", 404 => "0000000000000000", 405 => "0000000000000000", 406 => "0000000000000000", 407 => "0000000000000000", 408 => "0000000000000000", 409 => "0000000000000000", 410 => "0000000000000000", 411 => "0000000000000000", 412 => "0000000000000000", 413 => "0000000000000000", 414 => "0000000000000000", 415 => "0000000000000000", 416 => "0000000000000000", 417 => "0000000000000000", 418 => "0000000000000000", 419 => "0000000000000000", 420 => "0000000000000000", 421 => "0000000000000000", 422 => "0000000000000000", 423 => "0000000000000000", 424 => "0000000000000000", 425 => "0000000000000000", 426 => "0000000000000000", 427 => "0000000000000000", 428 => "0000000000000000", 429 => "0000000000000000", 430 => "0000000000000000", 431 => "0000000000000000", 432 => "0000000000000000", 433 => "0000000000000000", 434 => "0000000000000000", 435 => "0000000000000000", 436 => "0000000000000000", 437 => "0000000000000000", 438 => "0000000000000000", 439 => "0000000000000000", 440 => "0000000000000000", 441 => "0000000000000000", 442 => "0000000000000000", 443 => "0000000000000000", 444 => "0000000000000000", 445 => "0000000000000000", 446 => "0000000000000000", 447 => "0000000000000000", 448 => "0000000000000000", 449 => "0000000000000000", 450 => "0000000000000000", 451 => "0000000000000000", 452 => "0000000000000000", 453 => "0000000000000000", 454 => "0000000000000000", 455 => "0000000000000000", 456 => "0000000000000000", 457 => "0000000000000000", 458 => "0000000000000000", 459 => "0000000000000000", 460 => "0000000000000000", 461 => "0000000000000000", 462 => "0000000000000000", 463 => "0000000000000000", 464 => "0000000000000000", 465 => "0000000000000000", 466 => "0000000000000000", 467 => "0000000000000000", 468 => "0000000000000000", 469 => "0000000000000000", 470 => "0000000000000000", 471 => "0000000000000000", 472 => "0000000000000000", 473 => "0000000000000000", 474 => "0000000000000000", 475 => "0000000000000000", 476 => "0000000000000000", 477 => "0000000000000000", 478 => "0000000000000000", 479 => "0000000000000000", 480 => "0000000000000000", 481 => "0000000000000000", 482 => "0000000000000000", 483 => "0000000000000000", 484 => "0000000000000000", 485 => "0000000000000000", 486 => "0000000000000000", 487 => "0000000000000000", 488 => "0000000000000000", 489 => "0000000000000000", 490 => "0000000000000000", 491 => "0000000000000000", 492 => "0000000000000000", 493 => "0000000000000000", 494 => "0000000000000000", 495 => "0000000000000000", 496 => "0000000000000000", 497 => "0000000000000000", 498 => "0000000000000000", 499 => "0000000000000000", 500 => "0000000000000000", 501 => "0000000000000000", 502 => "0000000000000000", 503 => "0000000000000000", 504 => "0000000000000000", 505 => "0000000000000000", 506 => "0000000000000000", 507 => "0000000000000000", 508 => "0000000000000000", 509 => "0000000000000000", 510 => "0000000000000000", 511 => "0000000000000000", 512 => "0000000000000000", 513 => "0000000000000000", 514 => "0000000000000000", 515 => "0000000000000000", 516 => "0000000000000000", 517 => "0000000000000000", 518 => "0000000000000000", 519 => "0000000000000000", 520 => "0000000000000000", 521 => "0000000000000000", 522 => "0000000000000000", 523 => "0000000000000000", 524 => "0000000000000000", 525 => "0000000000000000", 526 => "0000000000000000", 527 => "0000000000000000", 528 => "0000000000000000", 529 => "0000000000000000", 530 => "0000000000000000", 531 => "0000000000000000", 532 => "0000000000000000", 533 => "0000000000000000", 534 => "0000000000000000", 535 => "0000000000000000", 536 => "0000000000000000", 537 => "0000000000000000", 538 => "0000000000000000", 539 => "0000000000000000", 540 => "0000000000000000", 541 => "0000000000000000", 542 => "0000000000000000", 543 => "0000000000000000", 544 => "0000000000000000", 545 => "0000000000000000", 546 => "0000000000000000", 547 => "0000000000000000", 548 => "0000000000000000", 549 => "0000000000000000", 550 => "0000000000000000", 551 => "0000000000000000", 552 => "0000000000000000", 553 => "0000000000000000", 554 => "0000000000000000", 555 => "0000000000000000", 556 => "0000000000000000", 557 => "0000000000000000", 558 => "0000000000000000", 559 => "0000000000000000", 560 => "0000000000000000", 561 => "0000000000000000", 562 => "0000000000000000", 563 => "0000000000000000", 564 => "0000000000000000", 565 => "0000000000000000", 566 => "0000000000000000", 567 => "0000000000000000", 568 => "0000000000000000", 569 => "0000000000000000", 570 => "0000000000000000", 571 => "0000000000000000", 572 => "0000000000000000", 573 => "0000000000000000", 574 => "0000000000000000", 575 => "0000000000000000", 576 => "0000000000000000", 577 => "0000000000000000", 578 => "0000000000000000", 579 => "0000000000000000", 580 => "0000000000000000", 581 => "0000000000000000", 582 => "0000000000000000", 583 => "0000000000000000", 584 => "0000000000000000", 585 => "0000000000000000", 586 => "0000000000000000", 587 => "0000000000000000", 588 => "0000000000000000", 589 => "0000000000000000", 590 => "0000000000000000", 591 => "0000000000000000", 592 => "0000000000000000", 593 => "0000000000000000", 594 => "0000000000000000", 595 => "0000000000000000", 596 => "0000000000000000", 597 => "0000000000000000", 598 => "0000000000000000", 599 => "0000000000000000", 600 => "0000000000000000", 601 => "0000000000000000", 602 => "0000000000000000", 603 => "0000000000000000", 604 => "0000000000000000", 605 => "0000000000000000", 606 => "0000000000000000", 607 => "0000000000000000", 608 => "0000000000000000", 609 => "0000000000000000", 610 => "0000000000000000", 611 => "0000000000000000", 612 => "0000000000000000", 613 => "0000000000000000", 614 => "0000000000000000", 615 => "0000000000000000", 616 => "0000000000000000", 617 => "0000000000000000", 618 => "0000000000000000", 619 => "0000000000000000", 620 => "0000000000000000", 621 => "0000000000000000", 622 => "0000000000000000", 623 => "0000000000000000", 624 => "0000000000000000", 625 => "0000000000000000", 626 => "0000000000000000", 627 => "0000000000000000", 628 => "0000000000000000", 629 => "0000000000000000", 630 => "0000000000000000", 631 => "0000000000000000", 632 => "0000000000000000", 633 => "0000000000000000", 634 => "0000000000000000", 635 => "0000000000000000", 636 => "0000000000000000", 637 => "0000000000000000", 638 => "0000000000000000", 639 => "0000000000000000", 640 => "0000000000000000", 641 => "0000000000000000", 642 => "0000000000000000", 643 => "0000000000000000", 644 => "0000000000000000", 645 => "0000000000000000", 646 => "0000000000000000", 647 => "0000000000000000", 648 => "0000000000000000", 649 => "0000000000000000", 650 => "0000000000000000", 651 => "0000000000000000", 652 => "0000000000000000", 653 => "0000000000000000", 654 => "0000000000000000", 655 => "0000000000000000", 656 => "0000000000000000", 657 => "0000000000000000", 658 => "0000000000000000", 659 => "0000000000000000", 660 => "0000000000000000", 661 => "0000000000000000", 662 => "0000000000000000", 663 => "0000000000000000", 664 => "0000000000000000", 665 => "0000000000000000", 666 => "0000000000000000", 667 => "0000000000000000", 668 => "0000000000000000", 669 => "0000000000000000", 670 => "0000000000000000", 671 => "0000000000000000", 672 => "0000000000000000", 673 => "0000000000000000", 674 => "0000000000000000", 675 => "0000000000000000", 676 => "0000000000000000", 677 => "0000000000000000", 678 => "0000000000000000", 679 => "0000000000000000", 680 => "0000000000000000", 681 => "0000000000000000", 682 => "0000000000000000", 683 => "0000000000000000", 684 => "0000000000000000", 685 => "0000000000000000", 686 => "0000000000000000", 687 => "0000000000000000", 688 => "0000000000000000", 689 => "0000000000000000", 690 => "0000000000000000", 691 => "0000000000000000", 692 => "0000000000000000", 693 => "0000000000000000", 694 => "0000000000000000", 695 => "0000000000000000", 696 => "0000000000000000", 697 => "0000000000000000", 698 => "0000000000000000", 699 => "0000000000000000", 700 => "0000000000000000", 701 => "0000000000000000", 702 => "0000000000000000", 703 => "0000000000000000", 704 => "0000000000000000", 705 => "0000000000000000", 706 => "0000000000000000", 707 => "0000000000000000", 708 => "0000000000000000", 709 => "0000000000000000", 710 => "0000000000000000", 711 => "0000000000000000", 712 => "0000000000000000", 713 => "0000000000000000", 714 => "0000000000000000", 715 => "0000000000000000", 716 => "0000000000000000", 717 => "0000000000000000", 718 => "0000000000000000", 719 => "0000000000000000", 720 => "0000000000000000", 721 => "0000000000000000", 722 => "0000000000000000", 723 => "0000000000000000", 724 => "0000000000000000", 725 => "0000000000000000", 726 => "0000000000000000", 727 => "0000000000000000", 728 => "0000000000000000", 729 => "0000000000000000", 730 => "0000000000000000", 731 => "0000000000000000", 732 => "0000000000000000", 733 => "0000000000000000", 734 => "0000000000000000", 735 => "0000000000000000", 736 => "0000000000000000", 737 => "0000000000000000", 738 => "0000000000000000", 739 => "0000000000000000", 740 => "0000000000000000", 741 => "0000000000000000", 742 => "0000000000000000", 743 => "0000000000000000", 744 => "0000000000000000", 745 => "0000000000000000", 746 => "0000000000000000", 747 => "0000000000000000", 748 => "0000000000000000", 749 => "0000000000000000", 750 => "0000000000000000", 751 => "0000000000000000", 752 => "0000000000000000", 753 => "0000000000000000", 754 => "0000000000000000", 755 => "0000000000000000", 756 => "0000000000000000", 757 => "0000000000000000", 758 => "0000000000000000", 759 => "0000000000000000", 760 => "0000000000000000", 761 => "0000000000000000", 762 => "0000000000000000", 763 => "0000000000000000", 764 => "0000000000000000", 765 => "0000000000000000", 766 => "0000000000000000", 767 => "0000000000000000", 768 => "0000000000000000", 769 => "0000000000000000", 770 => "0000000000000000", 771 => "0000000000000000", 772 => "0000000000000000", 773 => "0000000000000000", 774 => "0000000000000000", 775 => "0000000000000000", 776 => "0000000000000000", 777 => "0000000000000000", 778 => "0000000000000000", 779 => "0000000000000000", 780 => "0000000000000000", 781 => "0000000000000000", 782 => "0000000000000000", 783 => "0000000000000000", 784 => "0000000000000000", 785 => "0000000000000000", 786 => "0000000000000000", 787 => "0000000000000000", 788 => "0000000000000000", 789 => "0000000000000000", 790 => "0000000000000000", 791 => "0000000000000000", 792 => "0000000000000000", 793 => "0000000000000000", 794 => "0000000000000000", 795 => "0000000000000000", 796 => "0000000000000000", 797 => "0000000000000000", 798 => "0000000000000000", 799 => "0000000000000000", 800 => "0000000000000000", 801 => "0000000000000000", 802 => "0000000000000000", 803 => "0000000000000000", 804 => "0000000000000000", 805 => "0000000000000000", 806 => "0000000000000000", 807 => "0000000000000000", 808 => "0000000000000000", 809 => "0000000000000000", 810 => "0000000000000000", 811 => "0000000000000000", 812 => "0000000000000000", 813 => "0000000000000000", 814 => "0000000000000000", 815 => "0000000000000000", 816 => "0000000000000000", 817 => "0000000000000000", 818 => "0000000000000000", 819 => "0000000000000000", 820 => "0000000000000000", 821 => "0000000000000000", 822 => "0000000000000000", 823 => "0000000000000000", 824 => "0000000000000000", 825 => "0000000000000000", 826 => "0000000000000000", 827 => "0000000000000000", 828 => "0000000000000000", 829 => "0000000000000000", 830 => "0000000000000000", 831 => "0000000000000000", 832 => "0000000000000000", 833 => "0000000000000000", 834 => "0000000000000000", 835 => "0000000000000000", 836 => "0000000000000000", 837 => "0000000000000000", 838 => "0000000000000000", 839 => "0000000000000000", 840 => "0000000000000000", 841 => "0000000000000000", 842 => "0000000000000000", 843 => "0000000000000000", 844 => "0000000000000000", 845 => "0000000000000000", 846 => "0000000000000000", 847 => "0000000000000000", 848 => "0000000000000000", 849 => "0000000000000000", 850 => "0000000000000000", 851 => "0000000000000000", 852 => "0000000000000000", 853 => "0000000000000000", 854 => "0000000000000000", 855 => "0000000000000000", 856 => "0000000000000000", 857 => "0000000000000000", 858 => "0000000000000000", 859 => "0000000000000000", 860 => "0000000000000000", 861 => "0000000000000000", 862 => "0000000000000000", 863 => "0000000000000000", 864 => "0000000000000000", 865 => "0000000000000000", 866 => "0000000000000000", 867 => "0000000000000000", 868 => "0000000000000000", 869 => "0000000000000000", 870 => "0000000000000000", 871 => "0000000000000000", 872 => "0000000000000000", 873 => "0000000000000000", 874 => "0000000000000000", 875 => "0000000000000000", 876 => "0000000000000000", 877 => "0000000000000000", 878 => "0000000000000000", 879 => "0000000000000000", 880 => "0000000000000000", 881 => "0000000000000000", 882 => "0000000000000000", 883 => "0000000000000000", 884 => "0000000000000000", 885 => "0000000000000000", 886 => "0000000000000000", 887 => "0000000000000000", 888 => "0000000000000000", 889 => "0000000000000000", 890 => "0000000000000000", 891 => "0000000000000000", 892 => "0000000000000000", 893 => "0000000000000000", 894 => "0000000000000000", 895 => "0000000000000000", 896 => "0000000000000000", 897 => "0000000000000000", 898 => "0000000000000000", 899 => "0000000000000000", 900 => "0000000000000000", 901 => "0000000000000000", 902 => "0000000000000000", 903 => "0000000000000000", 904 => "0000000000000000", 905 => "0000000000000000", 906 => "0000000000000000", 907 => "0000000000000000", 908 => "0000000000000000", 909 => "0000000000000000", 910 => "0000000000000000", 911 => "0000000000000000", 912 => "0000000000000000", 913 => "0000000000000000", 914 => "0000000000000000", 915 => "0000000000000000", 916 => "0000000000000000", 917 => "0000000000000000", 918 => "0000000000000000", 919 => "0000000000000000", 920 => "0000000000000000", 921 => "0000000000000000", 922 => "0000000000000000", 923 => "0000000000000000", 924 => "0000000000000000", 925 => "0000000000000000", 926 => "0000000000000000", 927 => "0000000000000000", 928 => "0000000000000000", 929 => "0000000000000000", 930 => "0000000000000000", 931 => "0000000000000000", 932 => "0000000000000000", 933 => "0000000000000000", 934 => "0000000000000000", 935 => "0000000000000000", 936 => "0000000000000000", 937 => "0000000000000000", 938 => "0000000000000000", 939 => "0000000000000000", 940 => "0000000000000000", 941 => "0000000000000000", 942 => "0000000000000000", 943 => "0000000000000000", 944 => "0000000000000000", 945 => "0000000000000000", 946 => "0000000000000000", 947 => "0000000000000000", 948 => "0000000000000000", 949 => "0000000000000000", 950 => "0000000000000000", 951 => "0000000000000000", 952 => "0000000000000000", 953 => "0000000000000000", 954 => "0000000000000000", 955 => "0000000000000000", 956 => "0000000000000000", 957 => "0000000000000000", 958 => "0000000000000000", 959 => "0000000000000000", 960 => "0000000000000000", 961 => "0000000000000000", 962 => "0000000000000000", 963 => "0000000000000000", 964 => "0000000000000000", 965 => "0000000000000000", 966 => "0000000000000000", 967 => "0000000000000000", 968 => "0000000000000000", 969 => "0000000000000000", 970 => "0000000000000000", 971 => "0000000000000000", 972 => "0000000000000000", 973 => "0000000000000000", 974 => "0000000000000000", 975 => "0000000000000000", 976 => "0000000000000000", 977 => "0000000000000000", 978 => "0000000000000000", 979 => "0000000000000000", 980 => "0000000000000000", 981 => "0000000000000000", 982 => "0000000000000000", 983 => "0000000000000000", 984 => "0000000000000000", 985 => "0000000000000000", 986 => "0000000000000000", 987 => "0000000000000000", 988 => "0000000000000000", 989 => "0000000000000000", 990 => "0000000000000000", 991 => "0000000000000000", 992 => "0000000000000000", 993 => "0000000000000000", 994 => "0000000000000000", 995 => "0000000000000000", 996 => "0000000000000000", 997 => "0000000000000000", 998 => "0000000000000000", 999 => "0000000000000000", 1000 => "0000000000000000", 1001 => "0000000000000000", 1002 => "0000000000000000", 1003 => "0000000000000000", 1004 => "0000000000000000", 1005 => "0000000000000000", 1006 => "0000000000000000", 1007 => "0000000000000000", 1008 => "0000000000000000", 1009 => "0000000000000000", 1010 => "0000000000000000", 1011 => "0000000000000000", 1012 => "0000000000000000", 1013 => "0000000000000000", 1014 => "0000000000000000", 1015 => "0000000000000000", 1016 => "0000000000000000", 1017 => "0000000000000000", 1018 => "0000000000000000", 1019 => "0000000000000000", 1020 => "0000000000000000", 1021 => "0000000000000000", 1022 => "0000000000000000", 1023 => "0000000000000000", 1024 => "0000000000000000", 1025 => "0000000000000000", 1026 => "0000000000000000", 1027 => "0000000000000000", 1028 => "0000000000000000", 1029 => "0000000000000000", 1030 => "0000000000000000", 1031 => "0000000000000000", 1032 => "0000000000000000", 1033 => "0000000000000000", 1034 => "0000000000000000", 1035 => "0000000000000000", 1036 => "0000000000000000", 1037 => "0000000000000000", 1038 => "0000000000000000", 1039 => "0000000000000000", 1040 => "0000000000000000", 1041 => "0000000000000000", 1042 => "0000000000000000", 1043 => "0000000000000000", 1044 => "0000000000000000", 1045 => "0000000000000000", 1046 => "0000000000000000", 1047 => "0000000000000000", 1048 => "0000000000000000", 1049 => "0000000000000000", 1050 => "0000000000000000", 1051 => "0000000000000000", 1052 => "0000000000000000", 1053 => "0000000000000000", 1054 => "0000000000000000", 1055 => "0000000000000000", 1056 => "0000000000000000", 1057 => "0000000000000000", 1058 => "0000000000000000", 1059 => "0000000000000000", 1060 => "0000000000000000", 1061 => "0000000000000000", 1062 => "0000000000000000", 1063 => "0000000000000000", 1064 => "0000000000000000", 1065 => "0000000000000000", 1066 => "0000000000000000", 1067 => "0000000000000000", 1068 => "0000000000000000", 1069 => "0000000000000000", 1070 => "0000000000000000", 1071 => "0000000000000000", 1072 => "0000000000000000", 1073 => "0000000000000000", 1074 => "0000000000000000", 1075 => "0000000000000000", 1076 => "0000000000000000", 1077 => "0000000000000000", 1078 => "0000000000000000", 1079 => "0000000000000000", 1080 => "0000000000000000", 1081 => "0000000000000000", 1082 => "0000000000000000", 1083 => "0000000000000000", 1084 => "0000000000000000", 1085 => "0000000000000000", 1086 => "0000000000000000", 1087 => "0000000000000000", 1088 => "0000000000000000", 1089 => "0000000000000000", 1090 => "0000000000000000", 1091 => "0000000000000000", 1092 => "0000000000000000", 1093 => "0000000000000000", 1094 => "0000000000000000", 1095 => "0000000000000000", 1096 => "0000000000000000", 1097 => "0000000000000000", 1098 => "0000000000000000", 1099 => "0000000000000000", 1100 => "0000000000000000", 1101 => "0000000000000000", 1102 => "0000000000000000", 1103 => "0000000000000000", 1104 => "0000000000000000", 1105 => "0000000000000000", 1106 => "0000000000000000", 1107 => "0000000000000000", 1108 => "0000000000000000", 1109 => "0000000000000000", 1110 => "0000000000000000", 1111 => "0000000000000000", 1112 => "0000000000000000", 1113 => "0000000000000000", 1114 => "0000000000000000", 1115 => "0000000000000000", 1116 => "0000000000000000", 1117 => "0000000000000000", 1118 => "0000000000000000", 1119 => "0000000000000000", 1120 => "0000000000000000", 1121 => "0000000000000000", 1122 => "0000000000000000", 1123 => "0000000000000000", 1124 => "0000000000000000", 1125 => "0000000000000000", 1126 => "0000000000000000", 1127 => "0000000000000000", 1128 => "0000000000000000", 1129 => "0000000000000000", 1130 => "0000000000000000", 1131 => "0000000000000000", 1132 => "0000000000000000", 1133 => "0000000000000000", 1134 => "0000000000000000", 1135 => "0000000000000000", 1136 => "0000000000000000", 1137 => "0000000000000000", 1138 => "0000000000000000", 1139 => "0000000000000000", 1140 => "0000000000000000", 1141 => "0000000000000000", 1142 => "0000000000000000", 1143 => "0000000000000000", 1144 => "0000000000000000", 1145 => "0000000000000000", 1146 => "0000000000000000", 1147 => "0000000000000000", 1148 => "0000000000000000", 1149 => "0000000000000000", 1150 => "0000000000000000", 1151 => "0000000000000000", 1152 => "0000000000000000", 1153 => "0000000000000000", 1154 => "0000000000000000", 1155 => "0000000000000000", 1156 => "0000000000000000", 1157 => "0000000000000000", 1158 => "0000000000000000", 1159 => "0000000000000000", 1160 => "0000000000000000", 1161 => "0000000000000000", 1162 => "0000000000000000", 1163 => "0000000000000000", 1164 => "0000000000000000", 1165 => "0000000000000000", 1166 => "0000000000000000", 1167 => "0000000000000000", 1168 => "0000000000000000", 1169 => "0000000000000000", 1170 => "0000000000000000", 1171 => "0000000000000000", 1172 => "0000000000000000", 1173 => "0000000000000000", 1174 => "0000000000000000", 1175 => "0000000000000000", 1176 => "0000000000000000", 1177 => "0000000000000000", 1178 => "0000000000000000", 1179 => "0000000000000000", 1180 => "0000000000000000", 1181 => "0000000000000000", 1182 => "0000000000000000", 1183 => "0000000000000000", 1184 => "0000000000000000", 1185 => "0000000000000000", 1186 => "0000000000000000", 1187 => "0000000000000000", 1188 => "0000000000000000", 1189 => "0000000000000000", 1190 => "0000000000000000", 1191 => "0000000000000000", 1192 => "0000000000000000", 1193 => "0000000000000000", 1194 => "0000000000000000", 1195 => "0000000000000000", 1196 => "0000000000000000", 1197 => "0000000000000000", 1198 => "0000000000000000", 1199 => "0000000000000000", 1200 => "0000000000000000", 1201 => "0000000000000000", 1202 => "0000000000000000", 1203 => "0000000000000000", 1204 => "0000000000000000", 1205 => "0000000000000000", 1206 => "0000000000000000", 1207 => "0000000000000000", 1208 => "0000000000000000", 1209 => "0000000000000000", 1210 => "0000000000000000", 1211 => "0000000000000000", 1212 => "0000000000000000", 1213 => "0000000000000000", 1214 => "0000000000000000", 1215 => "0000000000000000", 1216 => "0000000000000000", 1217 => "0000000000000000", 1218 => "0000000000000000", 1219 => "0000000000000000", 1220 => "0000000000000000", 1221 => "0000000000000000", 1222 => "0000000000000000", 1223 => "0000000000000000", 1224 => "0000000000000000", 1225 => "0000000000000000", 1226 => "0000000000000000", 1227 => "0000000000000000", 1228 => "0000000000000000", 1229 => "0000000000000000", 1230 => "0000000000000000", 1231 => "0000000000000000", 1232 => "0000000000000000", 1233 => "0000000000000000", 1234 => "0000000000000000", 1235 => "0000000000000000", 1236 => "0000000000000000", 1237 => "0000000000000000", 1238 => "0000000000000000", 1239 => "0000000000000000", 1240 => "0000000000000000", 1241 => "0000000000000000", 1242 => "0000000000000000", 1243 => "0000000000000000", 1244 => "0000000000000000", 1245 => "0000000000000000", 1246 => "0000000000000000", 1247 => "0000000000000000", 1248 => "0000000000000000", 1249 => "0000000000000000", 1250 => "0000000000000000", 1251 => "0000000000000000", 1252 => "0000000000000000", 1253 => "0000000000000000", 1254 => "0000000000000000", 1255 => "0000000000000000", 1256 => "0000000000000000", 1257 => "0000000000000000", 1258 => "0000000000000000", 1259 => "0000000000000000", 1260 => "0000000000000000", 1261 => "0000000000000000", 1262 => "0000000000000000", 1263 => "0000000000000000", 1264 => "0000000000000000", 1265 => "0000000000000000", 1266 => "0000000000000000", 1267 => "0000000000000000", 1268 => "0000000000000000", 1269 => "0000000000000000", 1270 => "0000000000000000", 1271 => "0000000000000000", 1272 => "0000000000000000", 1273 => "0000000000000000", 1274 => "0000000000000000", 1275 => "0000000000000000", 1276 => "0000000000000000", 1277 => "0000000000000000", 1278 => "0000000000000000", 1279 => "0000000000000000", 1280 => "0000000000000000", 1281 => "0000000000000000", 1282 => "0000000000000000", 1283 => "0000000000000000", 1284 => "0000000000000000", 1285 => "0000000000000000", 1286 => "0000000000000000", 1287 => "0000000000000000", 1288 => "0000000000000000", 1289 => "0000000000000000", 1290 => "0000000000000000", 1291 => "0000000000000000", 1292 => "0000000000000000", 1293 => "0000000000000000", 1294 => "0000000000000000", 1295 => "0000000000000000", 1296 => "0000000000000000", 1297 => "0000000000000000", 1298 => "0000000000000000", 1299 => "0000000000000000", 1300 => "0000000000000000", 1301 => "0000000000000000", 1302 => "0000000000000000", 1303 => "0000000000000000", 1304 => "0000000000000000", 1305 => "0000000000000000", 1306 => "0000000000000000", 1307 => "0000000000000000", 1308 => "0000000000000000", 1309 => "0000000000000000", 1310 => "0000000000000000", 1311 => "0000000000000000", 1312 => "0000000000000000", 1313 => "0000000000000000", 1314 => "0000000000000000", 1315 => "0000000000000000", 1316 => "0000000000000000", 1317 => "0000000000000000", 1318 => "0000000000000000", 1319 => "0000000000000000", 1320 => "0000000000000000", 1321 => "0000000000000000", 1322 => "0000000000000000", 1323 => "0000000000000000", 1324 => "0000000000000000", 1325 => "0000000000000000", 1326 => "0000000000000000", 1327 => "0000000000000000", 1328 => "0000000000000000", 1329 => "0000000000000000", 1330 => "0000000000000000", 1331 => "0000000000000000", 1332 => "0000000000000000", 1333 => "0000000000000000", 1334 => "0000000000000000", 1335 => "0000000000000000", 1336 => "0000000000000000", 1337 => "0000000000000000", 1338 => "0000000000000000", 1339 => "0000000000000000", 1340 => "0000000000000000", 1341 => "0000000000000000", 1342 => "0000000000000000", 1343 => "0000000000000000", 1344 => "0000000000000000", 1345 => "0000000000000000", 1346 => "0000000000000000", 1347 => "0000000000000000", 1348 => "0000000000000000", 1349 => "0000000000000000", 1350 => "0000000000000000", 1351 => "0000000000000000", 1352 => "0000000000000000", 1353 => "0000000000000000", 1354 => "0000000000000000", 1355 => "0000000000000000", 1356 => "0000000000000000", 1357 => "0000000000000000", 1358 => "0000000000000000", 1359 => "0000000000000000", 1360 => "0000000000000000", 1361 => "0000000000000000", 1362 => "0000000000000000", 1363 => "0000000000000000", 1364 => "0000000000000000", 1365 => "0000000000000000", 1366 => "0000000000000000", 1367 => "0000000000000000", 1368 => "0000000000000000", 1369 => "0000000000000000", 1370 => "0000000000000000", 1371 => "0000000000000000", 1372 => "0000000000000000", 1373 => "0000000000000000", 1374 => "0000000000000000", 1375 => "0000000000000000", 1376 => "0000000000000000", 1377 => "0000000000000000", 1378 => "0000000000000000", 1379 => "0000000000000000", 1380 => "0000000000000000", 1381 => "0000000000000000", 1382 => "0000000000000000", 1383 => "0000000000000000", 1384 => "0000000000000000", 1385 => "0000000000000000", 1386 => "0000000000000000", 1387 => "0000000000000000", 1388 => "0000000000000000", 1389 => "0000000000000000", 1390 => "0000000000000000", 1391 => "0000000000000000", 1392 => "0000000000000000", 1393 => "0000000000000000", 1394 => "0000000000000000", 1395 => "0000000000000000", 1396 => "0000000000000000", 1397 => "0000000000000000", 1398 => "0000000000000000", 1399 => "0000000000000000", 1400 => "0000000000000000", 1401 => "0000000000000000", 1402 => "0000000000000000", 1403 => "0000000000000000", 1404 => "0000000000000000", 1405 => "0000000000000000", 1406 => "0000000000000000", 1407 => "0000000000000000", 1408 => "0000000000000000", 1409 => "0000000000000000", 1410 => "0000000000000000", 1411 => "0000000000000000", 1412 => "0000000000000000", 1413 => "0000000000000000", 1414 => "0000000000000000", 1415 => "0000000000000000", 1416 => "0000000000000000", 1417 => "0000000000000000", 1418 => "0000000000000000", 1419 => "0000000000000000", 1420 => "0000000000000000", 1421 => "0000000000000000", 1422 => "0000000000000000", 1423 => "0000000000000000", 1424 => "0000000000000000", 1425 => "0000000000000000", 1426 => "0000000000000000", 1427 => "0000000000000000", 1428 => "0000000000000000", 1429 => "0000000000000000", 1430 => "0000000000000000", 1431 => "0000000000000000", 1432 => "0000000000000000", 1433 => "0000000000000000", 1434 => "0000000000000000", 1435 => "0000000000000000", 1436 => "0000000000000000", 1437 => "0000000000000000", 1438 => "0000000000000000", 1439 => "0000000000000000", 1440 => "0000000000000000", 1441 => "0000000000000000", 1442 => "0000000000000000", 1443 => "0000000000000000", 1444 => "0000000000000000", 1445 => "0000000000000000", 1446 => "0000000000000000", 1447 => "0000000000000000", 1448 => "0000000000000000", 1449 => "0000000000000000", 1450 => "0000000000000000", 1451 => "0000000000000000", 1452 => "0000000000000000", 1453 => "0000000000000000", 1454 => "0000000000000000", 1455 => "0000000000000000", 1456 => "0000000000000000", 1457 => "0000000000000000", 1458 => "0000000000000000", 1459 => "0000000000000000", 1460 => "0000000000000000", 1461 => "0000000000000000", 1462 => "0000000000000000", 1463 => "0000000000000000", 1464 => "0000000000000000", 1465 => "0000000000000000", 1466 => "0000000000000000", 1467 => "0000000000000000", 1468 => "0000000000000000", 1469 => "0000000000000000", 1470 => "0000000000000000", 1471 => "0000000000000000", 1472 => "0000000000000000", 1473 => "0000000000000000", 1474 => "0000000000000000", 1475 => "0000000000000000", 1476 => "0000000000000000", 1477 => "0000000000000000", 1478 => "0000000000000000", 1479 => "0000000000000000", 1480 => "0000000000000000", 1481 => "0000000000000000", 1482 => "0000000000000000", 1483 => "0000000000000000", 1484 => "0000000000000000", 1485 => "0000000000000000", 1486 => "0000000000000000", 1487 => "0000000000000000", 1488 => "0000000000000000", 1489 => "0000000000000000", 1490 => "0000000000000000", 1491 => "0000000000000000", 1492 => "0000000000000000", 1493 => "0000000000000000", 1494 => "0000000000000000", 1495 => "0000000000000000", 1496 => "0000000000000000", 1497 => "0000000000000000", 1498 => "0000000000000000", 1499 => "0000000000000000", 1500 => "0000000000000000", 1501 => "0000000000000000", 1502 => "0000000000000000", 1503 => "0000000000000000", 1504 => "0000000000000000", 1505 => "0000000000000000", 1506 => "0000000000000000", 1507 => "0000000000000000", 1508 => "0000000000000000", 1509 => "0000000000000000", 1510 => "0000000000000000", 1511 => "0000000000000000", 1512 => "0000000000000000", 1513 => "0000000000000000", 1514 => "0000000000000000", 1515 => "0000000000000000", 1516 => "0000000000000000", 1517 => "0000000000000000", 1518 => "0000000000000000", 1519 => "0000000000000000", 1520 => "0000000000000000", 1521 => "0000000000000000", 1522 => "0000000000000000", 1523 => "0000000000000000", 1524 => "0000000000000000", 1525 => "0000000000000000", 1526 => "0000000000000000", 1527 => "0000000000000000", 1528 => "0000000000000000", 1529 => "0000000000000000", 1530 => "0000000000000000", 1531 => "0000000000000000", 1532 => "0000000000000000", 1533 => "0000000000000000", 1534 => "0000000000000000", 1535 => "0000000000000000", 1536 => "0000000000000000", 1537 => "0000000000000000", 1538 => "0000000000000000", 1539 => "0000000000000000", 1540 => "0000000000000000", 1541 => "0000000000000000", 1542 => "0000000000000000", 1543 => "0000000000000000", 1544 => "0000000000000000", 1545 => "0000000000000000", 1546 => "0000000000000000", 1547 => "0000000000000000", 1548 => "0000000000000000", 1549 => "0000000000000000", 1550 => "0000000000000000", 1551 => "0000000000000000", 1552 => "0000000000000000", 1553 => "0000000000000000", 1554 => "0000000000000000", 1555 => "0000000000000000", 1556 => "0000000000000000", 1557 => "0000000000000000", 1558 => "0000000000000000", 1559 => "0000000000000000", 1560 => "0000000000000000", 1561 => "0000000000000000", 1562 => "0000000000000000", 1563 => "0000000000000000", 1564 => "0000000000000000", 1565 => "0000000000000000", 1566 => "0000000000000000", 1567 => "0000000000000000", 1568 => "0000000000000000", 1569 => "0000000000000000", 1570 => "0000000000000000", 1571 => "0000000000000000", 1572 => "0000000000000000", 1573 => "0000000000000000", 1574 => "0000000000000000", 1575 => "0000000000000000", 1576 => "0000000000000000", 1577 => "0000000000000000", 1578 => "0000000000000000", 1579 => "0000000000000000", 1580 => "0000000000000000", 1581 => "0000000000000000", 1582 => "0000000000000000", 1583 => "0000000000000000", 1584 => "0000000000000000", 1585 => "0000000000000000", 1586 => "0000000000000000", 1587 => "0000000000000000", 1588 => "0000000000000000", 1589 => "0000000000000000", 1590 => "0000000000000000", 1591 => "0000000000000000", 1592 => "0000000000000000", 1593 => "0000000000000000", 1594 => "0000000000000000", 1595 => "0000000000000000", 1596 => "0000000000000000", 1597 => "0000000000000000", 1598 => "0000000000000000", 1599 => "0000000000000000", 1600 => "0000000000000000", 1601 => "0000000000000000", 1602 => "0000000000000000", 1603 => "0000000000000000", 1604 => "0000000000000000", 1605 => "0000000000000000", 1606 => "0000000000000000", 1607 => "0000000000000000", 1608 => "0000000000000000", 1609 => "0000000000000000", 1610 => "0000000000000000", 1611 => "0000000000000000", 1612 => "0000000000000000", 1613 => "0000000000000000", 1614 => "0000000000000000", 1615 => "0000000000000000", 1616 => "0000000000000000", 1617 => "0000000000000000", 1618 => "0000000000000000", 1619 => "0000000000000000", 1620 => "0000000000000000", 1621 => "0000000000000000", 1622 => "0000000000000000", 1623 => "0000000000000000", 1624 => "0000000000000000", 1625 => "0000000000000000", 1626 => "0000000000000000", 1627 => "0000000000000000", 1628 => "0000000000000000", 1629 => "0000000000000000", 1630 => "0000000000000000", 1631 => "0000000000000000", 1632 => "0000000000000000", 1633 => "0000000000000000", 1634 => "0000000000000000", 1635 => "0000000000000000", 1636 => "0000000000000000", 1637 => "0000000000000000", 1638 => "0000000000000000", 1639 => "0000000000000000", 1640 => "0000000000000000", 1641 => "0000000000000000", 1642 => "0000000000000000", 1643 => "0000000000000000", 1644 => "0000000000000000", 1645 => "0000000000000000", 1646 => "0000000000000000", 1647 => "0000000000000000", 1648 => "0000000000000000", 1649 => "0000000000000000", 1650 => "0000000000000000", 1651 => "0000000000000000", 1652 => "0000000000000000", 1653 => "0000000000000000", 1654 => "0000000000000000", 1655 => "0000000000000000", 1656 => "0000000000000000", 1657 => "0000000000000000", 1658 => "0000000000000000", 1659 => "0000000000000000", 1660 => "0000000000000000", 1661 => "0000000000000000", 1662 => "0000000000000000", 1663 => "0000000000000000", 1664 => "0000000000000000", 1665 => "0000000000000000", 1666 => "0000000000000000", 1667 => "0000000000000000", 1668 => "0000000000000000", 1669 => "0000000000000000", 1670 => "0000000000000000", 1671 => "0000000000000000", 1672 => "0000000000000000", 1673 => "0000000000000000", 1674 => "0000000000000000", 1675 => "0000000000000000", 1676 => "0000000000000000", 1677 => "0000000000000000", 1678 => "0000000000000000", 1679 => "0000000000000000", 1680 => "0000000000000000", 1681 => "0000000000000000", 1682 => "0000000000000000", 1683 => "0000000000000000", 1684 => "0000000000000000", 1685 => "0000000000000000", 1686 => "0000000000000000", 1687 => "0000000000000000", 1688 => "0000000000000000", 1689 => "0000000000000000", 1690 => "0000000000000000", 1691 => "0000000000000000", 1692 => "0000000000000000", 1693 => "0000000000000000", 1694 => "0000000000000000", 1695 => "0000000000000000", 1696 => "0000000000000000", 1697 => "0000000000000000", 1698 => "0000000000000000", 1699 => "0000000000000000", 1700 => "0000000000000000", 1701 => "0000000000000000", 1702 => "0000000000000000", 1703 => "0000000000000000", 1704 => "0000000000000000", 1705 => "0000000000000000", 1706 => "0000000000000000", 1707 => "0000000000000000", 1708 => "0000000000000000", 1709 => "0000000000000000", 1710 => "0000000000000000", 1711 => "0000000000000000", 1712 => "0000000000000000", 1713 => "0000000000000000", 1714 => "0000000000000000", 1715 => "0000000000000000", 1716 => "0000000000000000", 1717 => "0000000000000000", 1718 => "0000000000000000", 1719 => "0000000000000000", 1720 => "0000000000000000", 1721 => "0000000000000000", 1722 => "0000000000000000", 1723 => "0000000000000000", 1724 => "0000000000000000", 1725 => "0000000000000000", 1726 => "0000000000000000", 1727 => "0000000000000000", 1728 => "0000000000000000", 1729 => "0000000000000000", 1730 => "0000000000000000", 1731 => "0000000000000000", 1732 => "0000000000000000", 1733 => "0000000000000000", 1734 => "0000000000000000", 1735 => "0000000000000000", 1736 => "0000000000000000", 1737 => "0000000000000000", 1738 => "0000000000000000", 1739 => "0000000000000000", 1740 => "0000000000000000", 1741 => "0000000000000000", 1742 => "0000000000000000", 1743 => "0000000000000000", 1744 => "0000000000000000", 1745 => "0000000000000000", 1746 => "0000000000000000", 1747 => "0000000000000000", 1748 => "0000000000000000", 1749 => "0000000000000000", 1750 => "0000000000000000", 1751 => "0000000000000000", 1752 => "0000000000000000", 1753 => "0000000000000000", 1754 => "0000000000000000", 1755 => "0000000000000000", 1756 => "0000000000000000", 1757 => "0000000000000000", 1758 => "0000000000000000", 1759 => "0000000000000000", 1760 => "0000000000000000", 1761 => "0000000000000000", 1762 => "0000000000000000", 1763 => "0000000000000000", 1764 => "0000000000000000", 1765 => "0000000000000000", 1766 => "0000000000000000", 1767 => "0000000000000000", 1768 => "0000000000000000", 1769 => "0000000000000000", 1770 => "0000000000000000", 1771 => "0000000000000000", 1772 => "0000000000000000", 1773 => "0000000000000000", 1774 => "0000000000000000", 1775 => "0000000000000000", 1776 => "0000000000000000", 1777 => "0000000000000000", 1778 => "0000000000000000", 1779 => "0000000000000000", 1780 => "0000000000000000", 1781 => "0000000000000000", 1782 => "0000000000000000", 1783 => "0000000000000000", 1784 => "0000000000000000", 1785 => "0000000000000000", 1786 => "0000000000000000", 1787 => "0000000000000000", 1788 => "0000000000000000", 1789 => "0000000000000000", 1790 => "0000000000000000", 1791 => "0000000000000000", 1792 => "0000000000000000", 1793 => "0000000000000000", 1794 => "0000000000000000", 1795 => "0000000000000000", 1796 => "0000000000000000", 1797 => "0000000000000000", 1798 => "0000000000000000", 1799 => "0000000000000000", 1800 => "0000000000000000", 1801 => "0000000000000000", 1802 => "0000000000000000", 1803 => "0000000000000000", 1804 => "0000000000000000", 1805 => "0000000000000000", 1806 => "0000000000000000", 1807 => "0000000000000000", 1808 => "0000000000000000", 1809 => "0000000000000000", 1810 => "0000000000000000", 1811 => "0000000000000000", 1812 => "0000000000000000", 1813 => "0000000000000000", 1814 => "0000000000000000", 1815 => "0000000000000000", 1816 => "0000000000000000", 1817 => "0000000000000000", 1818 => "0000000000000000", 1819 => "0000000000000000", 1820 => "0000000000000000", 1821 => "0000000000000000", 1822 => "0000000000000000", 1823 => "0000000000000000", 1824 => "0000000000000000", 1825 => "0000000000000000", 1826 => "0000000000000000", 1827 => "0000000000000000", 1828 => "0000000000000000", 1829 => "0000000000000000", 1830 => "0000000000000000", 1831 => "0000000000000000", 1832 => "0000000000000000", 1833 => "0000000000000000", 1834 => "0000000000000000", 1835 => "0000000000000000", 1836 => "0000000000000000", 1837 => "0000000000000000", 1838 => "0000000000000000", 1839 => "0000000000000000", 1840 => "0000000000000000", 1841 => "0000000000000000", 1842 => "0000000000000000", 1843 => "0000000000000000", 1844 => "0000000000000000", 1845 => "0000000000000000", 1846 => "0000000000000000", 1847 => "0000000000000000", 1848 => "0000000000000000", 1849 => "0000000000000000", 1850 => "0000000000000000", 1851 => "0000000000000000", 1852 => "0000000000000000", 1853 => "0000000000000000", 1854 => "0000000000000000", 1855 => "0000000000000000", 1856 => "0000000000000000", 1857 => "0000000000000000", 1858 => "0000000000000000", 1859 => "0000000000000000", 1860 => "0000000000000000", 1861 => "0000000000000000", 1862 => "0000000000000000", 1863 => "0000000000000000", 1864 => "0000000000000000", 1865 => "0000000000000000", 1866 => "0000000000000000", 1867 => "0000000000000000", 1868 => "0000000000000000", 1869 => "0000000000000000", 1870 => "0000000000000000", 1871 => "0000000000000000", 1872 => "0000000000000000", 1873 => "0000000000000000", 1874 => "0000000000000000", 1875 => "0000000000000000", 1876 => "0000000000000000", 1877 => "0000000000000000", 1878 => "0000000000000000", 1879 => "0000000000000000", 1880 => "0000000000000000", 1881 => "0000000000000000", 1882 => "0000000000000000", 1883 => "0000000000000000", 1884 => "0000000000000000", 1885 => "0000000000000000", 1886 => "0000000000000000", 1887 => "0000000000000000", 1888 => "0000000000000000", 1889 => "0000000000000000", 1890 => "0000000000000000", 1891 => "0000000000000000", 1892 => "0000000000000000", 1893 => "0000000000000000", 1894 => "0000000000000000", 1895 => "0000000000000000", 1896 => "0000000000000000", 1897 => "0000000000000000", 1898 => "0000000000000000", 1899 => "0000000000000000", 1900 => "0000000000000000", 1901 => "0000000000000000", 1902 => "0000000000000000", 1903 => "0000000000000000", 1904 => "0000000000000000", 1905 => "0000000000000000", 1906 => "0000000000000000", 1907 => "0000000000000000", 1908 => "0000000000000000", 1909 => "0000000000000000", 1910 => "0000000000000000", 1911 => "0000000000000000", 1912 => "0000000000000000", 1913 => "0000000000000000", 1914 => "0000000000000000", 1915 => "0000000000000000", 1916 => "0000000000000000", 1917 => "0000000000000000", 1918 => "0000000000000000", 1919 => "0000000000000000", 1920 => "0000000000000000", 1921 => "0000000000000000", 1922 => "0000000000000000", 1923 => "0000000000000000", 1924 => "0000000000000000", 1925 => "0000000000000000", 1926 => "0000000000000000", 1927 => "0000000000000000", 1928 => "0000000000000000", 1929 => "0000000000000000", 1930 => "0000000000000000", 1931 => "0000000000000000", 1932 => "0000000000000000", 1933 => "0000000000000000", 1934 => "0000000000000000", 1935 => "0000000000000000", 1936 => "0000000000000000", 1937 => "0000000000000000", 1938 => "0000000000000000", 1939 => "0000000000000000", 1940 => "0000000000000000", 1941 => "0000000000000000", 1942 => "0000000000000000", 1943 => "0000000000000000", 1944 => "0000000000000000", 1945 => "0000000000000000", 1946 => "0000000000000000", 1947 => "0000000000000000", 1948 => "0000000000000000", 1949 => "0000000000000000", 1950 => "0000000000000000", 1951 => "0000000000000000", 1952 => "0000000000000000", 1953 => "0000000000000000", 1954 => "0000000000000000", 1955 => "0000000000000000", 1956 => "0000000000000000", 1957 => "0000000000000000", 1958 => "0000000000000000", 1959 => "0000000000000000", 1960 => "0000000000000000", 1961 => "0000000000000000", 1962 => "0000000000000000", 1963 => "0000000000000000", 1964 => "0000000000000000", 1965 => "0000000000000000", 1966 => "0000000000000000", 1967 => "0000000000000000", 1968 => "0000000000000000", 1969 => "0000000000000000", 1970 => "0000000000000000", 1971 => "0000000000000000", 1972 => "0000000000000000", 1973 => "0000000000000000", 1974 => "0000000000000000", 1975 => "0000000000000000", 1976 => "0000000000000000", 1977 => "0000000000000000", 1978 => "0000000000000000", 1979 => "0000000000000000", 1980 => "0000000000000000", 1981 => "0000000000000000", 1982 => "0000000000000000", 1983 => "0000000000000000", 1984 => "0000000000000000", 1985 => "0000000000000000", 1986 => "0000000000000000", 1987 => "0000000000000000", 1988 => "0000000000000000", 1989 => "0000000000000000", 1990 => "0000000000000000", 1991 => "0000000000000000", 1992 => "0000000000000000", 1993 => "0000000000000000", 1994 => "0000000000000000", 1995 => "0000000000000000", 1996 => "0000000000000000", 1997 => "0000000000000000", 1998 => "0000000000000000", 1999 => "0000000000000000", 2000 => "0000000000000000", 2001 => "0000000000000000", 2002 => "0000000000000000", 2003 => "0000000000000000", 2004 => "0000000000000000", 2005 => "0000000000000000", 2006 => "0000000000000000", 2007 => "0000000000000000", 2008 => "0000000000000000", 2009 => "0000000000000000", 2010 => "0000000000000000", 2011 => "0000000000000000", 2012 => "0000000000000000", 2013 => "0000000000000000", 2014 => "0000000000000000", 2015 => "0000000000000000", 2016 => "0000000000000000", 2017 => "0000000000000000", 2018 => "0000000000000000", 2019 => "0000000000000000", 2020 => "0000000000000000", 2021 => "0000000000000000", 2022 => "0000000000000000", 2023 => "0000000000000000", 2024 => "0000000000000000", 2025 => "0000000000000000", 2026 => "0000000000000000", 2027 => "0000000000000000", 2028 => "0000000000000000", 2029 => "0000000000000000", 2030 => "0000000000000000", 2031 => "0000000000000000", 2032 => "0000000000000000", 2033 => "0000000000000000", 2034 => "0000000000000000", 2035 => "0000000000000000", 2036 => "0000000000000000", 2037 => "0000000000000000", 2038 => "0000000000000000", 2039 => "0000000000000000", 2040 => "0000000000000000", 2041 => "0000000000000000", 2042 => "0000000000000000", 2043 => "0000000000000000", 2044 => "0000000000000000", 2045 => "0000000000000000", 2046 => "0000000000000000", 2047 => "0000000000000000", 2048 => "0000000000000000", 2049 => "0000000000000000", 2050 => "0000000000000000", 2051 => "0000000000000000", 2052 => "0000000000000000", 2053 => "0000000000000000", 2054 => "0000000000000000", 2055 => "0000000000000000", 2056 => "0000000000000000", 2057 => "0000000000000000", 2058 => "0000000000000000", 2059 => "0000000000000000", 2060 => "0000000000000000", 2061 => "0000000000000000", 2062 => "0000000000000000", 2063 => "0000000000000000", 2064 => "0000000000000000", 2065 => "0000000000000000", 2066 => "0000000000000000", 2067 => "0000000000000000", 2068 => "0000000000000000", 2069 => "0000000000000000", 2070 => "0000000000000000", 2071 => "0000000000000000", 2072 => "0000000000000000", 2073 => "0000000000000000", 2074 => "0000000000000000", 2075 => "0000000000000000", 2076 => "0000000000000000", 2077 => "0000000000000000", 2078 => "0000000000000000", 2079 => "0000000000000000", 2080 => "0000000000000000", 2081 => "0000000000000000", 2082 => "0000000000000000", 2083 => "0000000000000000", 2084 => "0000000000000000", 2085 => "0000000000000000", 2086 => "0000000000000000", 2087 => "0000000000000000", 2088 => "0000000000000000", 2089 => "0000000000000000", 2090 => "0000000000000000", 2091 => "0000000000000000", 2092 => "0000000000000000", 2093 => "0000000000000000", 2094 => "0000000000000000", 2095 => "0000000000000000", 2096 => "0000000000000000", 2097 => "0000000000000000", 2098 => "0000000000000000", 2099 => "0000000000000000", 2100 => "0000000000000000", 2101 => "0000000000000000", 2102 => "0000000000000000", 2103 => "0000000000000000", 2104 => "0000000000000000", 2105 => "0000000000000000", 2106 => "0000000000000000", 2107 => "0000000000000000", 2108 => "0000000000000000", 2109 => "0000000000000000", 2110 => "0000000000000000", 2111 => "0000000000000000", 2112 => "0000000000000000", 2113 => "0000000000000000", 2114 => "0000000000000000", 2115 => "0000000000000000", 2116 => "0000000000000000", 2117 => "0000000000000000", 2118 => "0000000000000000", 2119 => "0000000000000000", 2120 => "0000000000000000", 2121 => "0000000000000000", 2122 => "0000000000000000", 2123 => "0000000000000000", 2124 => "0000000000000000", 2125 => "0000000000000000", 2126 => "0000000000000000", 2127 => "0000000000000000", 2128 => "0000000000000000", 2129 => "0000000000000000", 2130 => "0000000000000000", 2131 => "0000000000000000", 2132 => "0000000000000000", 2133 => "0000000000000000", 2134 => "0000000000000000", 2135 => "0000000000000000", 2136 => "0000000000000000", 2137 => "0000000000000000", 2138 => "0000000000000000", 2139 => "0000000000000000", 2140 => "0000000000000000", 2141 => "0000000000000000", 2142 => "0000000000000000", 2143 => "0000000000000000", 2144 => "0000000000000000", 2145 => "0000000000000000", 2146 => "0000000000000000", 2147 => "0000000000000000", 2148 => "0000000000000000", 2149 => "0000000000000000", 2150 => "0000000000000000", 2151 => "0000000000000000", 2152 => "0000000000000000", 2153 => "0000000000000000", 2154 => "0000000000000000", 2155 => "0000000000000000", 2156 => "0000000000000000", 2157 => "0000000000000000", 2158 => "0000000000000000", 2159 => "0000000000000000", 2160 => "0000000000000000", 2161 => "0000000000000000", 2162 => "0000000000000000", 2163 => "0000000000000000", 2164 => "0000000000000000", 2165 => "0000000000000000", 2166 => "0000000000000000", 2167 => "0000000000000000", 2168 => "0000000000000000", 2169 => "0000000000000000", 2170 => "0000000000000000", 2171 => "0000000000000000", 2172 => "0000000000000000", 2173 => "0000000000000000", 2174 => "0000000000000000", 2175 => "0000000000000000", 2176 => "0000000000000000", 2177 => "0000000000000000", 2178 => "0000000000000000", 2179 => "0000000000000000", 2180 => "0000000000000000", 2181 => "0000000000000000", 2182 => "0000000000000000", 2183 => "0000000000000000", 2184 => "0000000000000000", 2185 => "0000000000000000", 2186 => "0000000000000000", 2187 => "0000000000000000", 2188 => "0000000000000000", 2189 => "0000000000000000", 2190 => "0000000000000000", 2191 => "0000000000000000", 2192 => "0000000000000000", 2193 => "0000000000000000", 2194 => "0000000000000000", 2195 => "0000000000000000", 2196 => "0000000000000000", 2197 => "0000000000000000", 2198 => "0000000000000000", 2199 => "0000000000000000", 2200 => "0000000000000000", 2201 => "0000000000000000", 2202 => "0000000000000000", 2203 => "0000000000000000", 2204 => "0000000000000000", 2205 => "0000000000000000", 2206 => "0000000000000000", 2207 => "0000000000000000", 2208 => "0000000000000000", 2209 => "0000000000000000", 2210 => "0000000000000000", 2211 => "0000000000000000", 2212 => "0000000000000000", 2213 => "0000000000000000", 2214 => "0000000000000000", 2215 => "0000000000000000", 2216 => "0000000000000000", 2217 => "0000000000000000", 2218 => "0000000000000000", 2219 => "0000000000000000", 2220 => "0000000000000000", 2221 => "0000000000000000", 2222 => "0000000000000000", 2223 => "0000000000000000", 2224 => "0000000000000000", 2225 => "0000000000000000", 2226 => "0000000000000000", 2227 => "0000000000000000", 2228 => "0000000000000000", 2229 => "0000000000000000", 2230 => "0000000000000000", 2231 => "0000000000000000", 2232 => "0000000000000000", 2233 => "0000000000000000", 2234 => "0000000000000000", 2235 => "0000000000000000", 2236 => "0000000000000000", 2237 => "0000000000000000", 2238 => "0000000000000000", 2239 => "0000000000000000", 2240 => "0000000000000000", 2241 => "0000000000000000", 2242 => "0000000000000000", 2243 => "0000000000000000", 2244 => "0000000000000000", 2245 => "0000000000000000", 2246 => "0000000000000000", 2247 => "0000000000000000", 2248 => "0000000000000000", 2249 => "0000000000000000", 2250 => "0000000000000000", 2251 => "0000000000000000", 2252 => "0000000000000000", 2253 => "0000000000000000", 2254 => "0000000000000000", 2255 => "0000000000000000", 2256 => "0000000000000000", 2257 => "0000000000000000", 2258 => "0000000000000000", 2259 => "0000000000000000", 2260 => "0000000000000000", 2261 => "0000000000000000", 2262 => "0000000000000000", 2263 => "0000000000000000", 2264 => "0000000000000000", 2265 => "0000000000000000", 2266 => "0000000000000000", 2267 => "0000000000000000", 2268 => "0000000000000000", 2269 => "0000000000000000", 2270 => "0000000000000000", 2271 => "0000000000000000", 2272 => "0000000000000000", 2273 => "0000000000000000", 2274 => "0000000000000000", 2275 => "0000000000000000", 2276 => "0000000000000000", 2277 => "0000000000000000", 2278 => "0000000000000000", 2279 => "0000000000000000", 2280 => "0000000000000000", 2281 => "0000000000000000", 2282 => "0000000000000000", 2283 => "0000000000000000", 2284 => "0000000000000000", 2285 => "0000000000000000", 2286 => "0000000000000000", 2287 => "0000000000000000", 2288 => "0000000000000000", 2289 => "0000000000000000", 2290 => "0000000000000000", 2291 => "0000000000000000", 2292 => "0000000000000000", 2293 => "0000000000000000", 2294 => "0000000000000000", 2295 => "0000000000000000", 2296 => "0000000000000000", 2297 => "0000000000000000", 2298 => "0000000000000000", 2299 => "0000000000000000", 2300 => "0000000000000000", 2301 => "0000000000000000", 2302 => "0000000000000000", 2303 => "0000000000000000", 2304 => "0000000000000000", 2305 => "0000000000000000", 2306 => "0000000000000000", 2307 => "0000000000000000", 2308 => "0000000000000000", 2309 => "0000000000000000", 2310 => "0000000000000000", 2311 => "0000000000000000", 2312 => "0000000000000000", 2313 => "0000000000000000", 2314 => "0000000000000000", 2315 => "0000000000000000", 2316 => "0000000000000000", 2317 => "0000000000000000", 2318 => "0000000000000000", 2319 => "0000000000000000", 2320 => "0000000000000000", 2321 => "0000000000000000", 2322 => "0000000000000000", 2323 => "0000000000000000", 2324 => "0000000000000000", 2325 => "0000000000000000", 2326 => "0000000000000000", 2327 => "0000000000000000", 2328 => "0000000000000000", 2329 => "0000000000000000", 2330 => "0000000000000000", 2331 => "0000000000000000", 2332 => "0000000000000000", 2333 => "0000000000000000", 2334 => "0000000000000000", 2335 => "0000000000000000", 2336 => "0000000000000000", 2337 => "0000000000000000", 2338 => "0000000000000000", 2339 => "0000000000000000", 2340 => "0000000000000000", 2341 => "0000000000000000", 2342 => "0000000000000000", 2343 => "0000000000000000", 2344 => "0000000000000000", 2345 => "0000000000000000", 2346 => "0000000000000000", 2347 => "0000000000000000", 2348 => "0000000000000000", 2349 => "0000000000000000", 2350 => "0000000000000000", 2351 => "0000000000000000", 2352 => "0000000000000000", 2353 => "0000000000000000", 2354 => "0000000000000000", 2355 => "0000000000000000", 2356 => "0000000000000000", 2357 => "0000000000000000", 2358 => "0000000000000000", 2359 => "0000000000000000", 2360 => "0000000000000000", 2361 => "0000000000000000", 2362 => "0000000000000000", 2363 => "0000000000000000", 2364 => "0000000000000000", 2365 => "0000000000000000", 2366 => "0000000000000000", 2367 => "0000000000000000", 2368 => "0000000000000000", 2369 => "0000000000000000", 2370 => "0000000000000000", 2371 => "0000000000000000", 2372 => "0000000000000000", 2373 => "0000000000000000", 2374 => "0000000000000000", 2375 => "0000000000000000", 2376 => "0000000000000000", 2377 => "0000000000000000", 2378 => "0000000000000000", 2379 => "0000000000000000", 2380 => "0000000000000000", 2381 => "0000000000000000", 2382 => "0000000000000000", 2383 => "0000000000000000", 2384 => "0000000000000000", 2385 => "0000000000000000", 2386 => "0000000000000000", 2387 => "0000000000000000", 2388 => "0000000000000000", 2389 => "0000000000000000", 2390 => "0000000000000000", 2391 => "0000000000000000", 2392 => "0000000000000000", 2393 => "0000000000000000", 2394 => "0000000000000000", 2395 => "0000000000000000", 2396 => "0000000000000000", 2397 => "0000000000000000", 2398 => "0000000000000000", 2399 => "0000000000000000", 2400 => "0000000000000000", 2401 => "0000000000000000", 2402 => "0000000000000000", 2403 => "0000000000000000", 2404 => "0000000000000000", 2405 => "0000000000000000", 2406 => "0000000000000000", 2407 => "0000000000000000", 2408 => "0000000000000000", 2409 => "0000000000000000", 2410 => "0000000000000000", 2411 => "0000000000000000", 2412 => "0000000000000000", 2413 => "0000000000000000", 2414 => "0000000000000000", 2415 => "0000000000000000", 2416 => "0000000000000000", 2417 => "0000000000000000", 2418 => "0000000000000000", 2419 => "0000000000000000", 2420 => "0000000000000000", 2421 => "0000000000000000", 2422 => "0000000000000000", 2423 => "0000000000000000", 2424 => "0000000000000000", 2425 => "0000000000000000", 2426 => "0000000000000000", 2427 => "0000000000000000", 2428 => "0000000000000000", 2429 => "0000000000000000", 2430 => "0000000000000000", 2431 => "0000000000000000", 2432 => "0000000000000000", 2433 => "0000000000000000", 2434 => "0000000000000000", 2435 => "0000000000000000", 2436 => "0000000000000000", 2437 => "0000000000000000", 2438 => "0000000000000000", 2439 => "0000000000000000", 2440 => "0000000000000000", 2441 => "0000000000000000", 2442 => "0000000000000000", 2443 => "0000000000000000", 2444 => "0000000000000000", 2445 => "0000000000000000", 2446 => "0000000000000000", 2447 => "0000000000000000", 2448 => "0000000000000000", 2449 => "0000000000000000", 2450 => "0000000000000000", 2451 => "0000000000000000", 2452 => "0000000000000000", 2453 => "0000000000000000", 2454 => "0000000000000000", 2455 => "0000000000000000", 2456 => "0000000000000000", 2457 => "0000000000000000", 2458 => "0000000000000000", 2459 => "0000000000000000", 2460 => "0000000000000000", 2461 => "0000000000000000", 2462 => "0000000000000000", 2463 => "0000000000000000", 2464 => "0000000000000000", 2465 => "0000000000000000", 2466 => "0000000000000000", 2467 => "0000000000000000", 2468 => "0000000000000000", 2469 => "0000000000000000", 2470 => "0000000000000000", 2471 => "0000000000000000", 2472 => "0000000000000000", 2473 => "0000000000000000", 2474 => "0000000000000000", 2475 => "0000000000000000", 2476 => "0000000000000000", 2477 => "0000000000000000", 2478 => "0000000000000000", 2479 => "0000000000000000", 2480 => "0000000000000000", 2481 => "0000000000000000", 2482 => "0000000000000000", 2483 => "0000000000000000", 2484 => "0000000000000000", 2485 => "0000000000000000", 2486 => "0000000000000000", 2487 => "0000000000000000", 2488 => "0000000000000000", 2489 => "0000000000000000", 2490 => "0000000000000000", 2491 => "0000000000000000", 2492 => "0000000000000000", 2493 => "0000000000000000", 2494 => "0000000000000000", 2495 => "0000000000000000", 2496 => "0000000000000000", 2497 => "0000000000000000", 2498 => "0000000000000000", 2499 => "0000000000000000", 2500 => "0000000000000000", 2501 => "0000000000000000", 2502 => "0000000000000000", 2503 => "0000000000000000", 2504 => "0000000000000000", 2505 => "0000000000000000", 2506 => "0000000000000000", 2507 => "0000000000000000", 2508 => "0000000000000000", 2509 => "0000000000000000", 2510 => "0000000000000000", 2511 => "0000000000000000", 2512 => "0000000000000000", 2513 => "0000000000000000", 2514 => "0000000000000000", 2515 => "0000000000000000", 2516 => "0000000000000000", 2517 => "0000000000000000", 2518 => "0000000000000000", 2519 => "0000000000000000", 2520 => "0000000000000000", 2521 => "0000000000000000", 2522 => "0000000000000000", 2523 => "0000000000000000", 2524 => "0000000000000000", 2525 => "0000000000000000", 2526 => "0000000000000000", 2527 => "0000000000000000", 2528 => "0000000000000000", 2529 => "0000000000000000", 2530 => "0000000000000000", 2531 => "0000000000000000", 2532 => "0000000000000000", 2533 => "0000000000000000", 2534 => "0000000000000000", 2535 => "0000000000000000", 2536 => "0000000000000000", 2537 => "0000000000000000", 2538 => "0000000000000000", 2539 => "0000000000000000", 2540 => "0000000000000000", 2541 => "0000000000000000", 2542 => "0000000000000000", 2543 => "0000000000000000", 2544 => "0000000000000000", 2545 => "0000000000000000", 2546 => "0000000000000000", 2547 => "0000000000000000", 2548 => "0000000000000000", 2549 => "0000000000000000", 2550 => "0000000000000000", 2551 => "0000000000000000", 2552 => "0000000000000000", 2553 => "0000000000000000", 2554 => "0000000000000000", 2555 => "0000000000000000", 2556 => "0000000000000000", 2557 => "0000000000000000", 2558 => "0000000000000000", 2559 => "0000000000000000", 2560 => "0000000000000000", 2561 => "0000000000000000", 2562 => "0000000000000000", 2563 => "0000000000000000", 2564 => "0000000000000000", 2565 => "0000000000000000", 2566 => "0000000000000000", 2567 => "0000000000000000", 2568 => "0000000000000000", 2569 => "0000000000000000", 2570 => "0000000000000000", 2571 => "0000000000000000", 2572 => "0000000000000000", 2573 => "0000000000000000", 2574 => "0000000000000000", 2575 => "0000000000000000", 2576 => "0000000000000000", 2577 => "0000000000000000", 2578 => "0000000000000000", 2579 => "0000000000000000", 2580 => "0000000000000000", 2581 => "0000000000000000", 2582 => "0000000000000000", 2583 => "0000000000000000", 2584 => "0000000000000000", 2585 => "0000000000000000", 2586 => "0000000000000000", 2587 => "0000000000000000", 2588 => "0000000000000000", 2589 => "0000000000000000", 2590 => "0000000000000000", 2591 => "0000000000000000", 2592 => "0000000000000000", 2593 => "0000000000000000", 2594 => "0000000000000000", 2595 => "0000000000000000", 2596 => "0000000000000000", 2597 => "0000000000000000", 2598 => "0000000000000000", 2599 => "0000000000000000", 2600 => "0000000000000000", 2601 => "0000000000000000", 2602 => "0000000000000000", 2603 => "0000000000000000", 2604 => "0000000000000000", 2605 => "0000000000000000", 2606 => "0000000000000000", 2607 => "0000000000000000", 2608 => "0000000000000000", 2609 => "0000000000000000", 2610 => "0000000000000000", 2611 => "0000000000000000", 2612 => "0000000000000000", 2613 => "0000000000000000", 2614 => "0000000000000000", 2615 => "0000000000000000", 2616 => "0000000000000000", 2617 => "0000000000000000", 2618 => "0000000000000000", 2619 => "0000000000000000", 2620 => "0000000000000000", 2621 => "0000000000000000", 2622 => "0000000000000000", 2623 => "0000000000000000", 2624 => "0000000000000000", 2625 => "0000000000000000", 2626 => "0000000000000000", 2627 => "0000000000000000", 2628 => "0000000000000000", 2629 => "0000000000000000", 2630 => "0000000000000000", 2631 => "0000000000000000", 2632 => "0000000000000000", 2633 => "0000000000000000", 2634 => "0000000000000000", 2635 => "0000000000000000", 2636 => "0000000000000000", 2637 => "0000000000000000", 2638 => "0000000000000000", 2639 => "0000000000000000", 2640 => "0000000000000000", 2641 => "0000000000000000", 2642 => "0000000000000000", 2643 => "0000000000000000", 2644 => "0000000000000000", 2645 => "0000000000000000", 2646 => "0000000000000000", 2647 => "0000000000000000", 2648 => "0000000000000000", 2649 => "0000000000000000", 2650 => "0000000000000000", 2651 => "0000000000000000", 2652 => "0000000000000000", 2653 => "0000000000000000", 2654 => "0000000000000000", 2655 => "0000000000000000", 2656 => "0000000000000000", 2657 => "0000000000000000", 2658 => "0000000000000000", 2659 => "0000000000000000", 2660 => "0000000000000000", 2661 => "0000000000000000", 2662 => "0000000000000000", 2663 => "0000000000000000", 2664 => "0000000000000000", 2665 => "0000000000000000", 2666 => "0000000000000000", 2667 => "0000000000000000", 2668 => "0000000000000000", 2669 => "0000000000000000", 2670 => "0000000000000000", 2671 => "0000000000000000", 2672 => "0000000000000000", 2673 => "0000000000000000", 2674 => "0000000000000000", 2675 => "0000000000000000", 2676 => "0000000000000000", 2677 => "0000000000000000", 2678 => "0000000000000000", 2679 => "0000000000000000", 2680 => "0000000000000000", 2681 => "0000000000000000", 2682 => "0000000000000000", 2683 => "0000000000000000", 2684 => "0000000000000000", 2685 => "0000000000000000", 2686 => "0000000000000000", 2687 => "0000000000000000", 2688 => "0000000000000000", 2689 => "0000000000000000", 2690 => "0000000000000000", 2691 => "0000000000000000", 2692 => "0000000000000000", 2693 => "0000000000000000", 2694 => "0000000000000000", 2695 => "0000000000000000", 2696 => "0000000000000000", 2697 => "0000000000000000", 2698 => "0000000000000000", 2699 => "0000000000000000", 2700 => "0000000000000000", 2701 => "0000000000000000", 2702 => "0000000000000000", 2703 => "0000000000000000", 2704 => "0000000000000000", 2705 => "0000000000000000", 2706 => "0000000000000000", 2707 => "0000000000000000", 2708 => "0000000000000000", 2709 => "0000000000000000", 2710 => "0000000000000000", 2711 => "0000000000000000", 2712 => "0000000000000000", 2713 => "0000000000000000", 2714 => "0000000000000000", 2715 => "0000000000000000", 2716 => "0000000000000000", 2717 => "0000000000000000", 2718 => "0000000000000000", 2719 => "0000000000000000", 2720 => "0000000000000000", 2721 => "0000000000000000", 2722 => "0000000000000000", 2723 => "0000000000000000", 2724 => "0000000000000000", 2725 => "0000000000000000", 2726 => "0000000000000000", 2727 => "0000000000000000", 2728 => "0000000000000000", 2729 => "0000000000000000", 2730 => "0000000000000000", 2731 => "0000000000000000", 2732 => "0000000000000000", 2733 => "0000000000000000", 2734 => "0000000000000000", 2735 => "0000000000000000", 2736 => "0000000000000000", 2737 => "0000000000000000", 2738 => "0000000000000000", 2739 => "0000000000000000", 2740 => "0000000000000000", 2741 => "0000000000000000", 2742 => "0000000000000000", 2743 => "0000000000000000", 2744 => "0000000000000000", 2745 => "0000000000000000", 2746 => "0000000000000000", 2747 => "0000000000000000", 2748 => "0000000000000000", 2749 => "0000000000000000", 2750 => "0000000000000000", 2751 => "0000000000000000", 2752 => "0000000000000000", 2753 => "0000000000000000", 2754 => "0000000000000000", 2755 => "0000000000000000", 2756 => "0000000000000000", 2757 => "0000000000000000", 2758 => "0000000000000000", 2759 => "0000000000000000", 2760 => "0000000000000000", 2761 => "0000000000000000", 2762 => "0000000000000000", 2763 => "0000000000000000", 2764 => "0000000000000000", 2765 => "0000000000000000", 2766 => "0000000000000000", 2767 => "0000000000000000", 2768 => "0000000000000000", 2769 => "0000000000000000", 2770 => "0000000000000000", 2771 => "0000000000000000", 2772 => "0000000000000000", 2773 => "0000000000000000", 2774 => "0000000000000000", 2775 => "0000000000000000", 2776 => "0000000000000000", 2777 => "0000000000000000", 2778 => "0000000000000000", 2779 => "0000000000000000", 2780 => "0000000000000000", 2781 => "0000000000000000", 2782 => "0000000000000000", 2783 => "0000000000000000", 2784 => "0000000000000000", 2785 => "0000000000000000", 2786 => "0000000000000000", 2787 => "0000000000000000", 2788 => "0000000000000000", 2789 => "0000000000000000", 2790 => "0000000000000000", 2791 => "0000000000000000", 2792 => "0000000000000000", 2793 => "0000000000000000", 2794 => "0000000000000000", 2795 => "0000000000000000", 2796 => "0000000000000000", 2797 => "0000000000000000", 2798 => "0000000000000000", 2799 => "0000000000000000", 2800 => "0000000000000000", 2801 => "0000000000000000", 2802 => "0000000000000000", 2803 => "0000000000000000", 2804 => "0000000000000000", 2805 => "0000000000000000", 2806 => "0000000000000000", 2807 => "0000000000000000", 2808 => "0000000000000000", 2809 => "0000000000000000", 2810 => "0000000000000000", 2811 => "0000000000000000", 2812 => "0000000000000000", 2813 => "0000000000000000", 2814 => "0000000000000000", 2815 => "0000000000000000", 2816 => "0000000000000000", 2817 => "0000000000000000", 2818 => "0000000000000000", 2819 => "0000000000000000", 2820 => "0000000000000000", 2821 => "0000000000000000", 2822 => "0000000000000000", 2823 => "0000000000000000", 2824 => "0000000000000000", 2825 => "0000000000000000", 2826 => "0000000000000000", 2827 => "0000000000000000", 2828 => "0000000000000000", 2829 => "0000000000000000", 2830 => "0000000000000000", 2831 => "0000000000000000", 2832 => "0000000000000000", 2833 => "0000000000000000", 2834 => "0000000000000000", 2835 => "0000000000000000", 2836 => "0000000000000000", 2837 => "0000000000000000", 2838 => "0000000000000000", 2839 => "0000000000000000", 2840 => "0000000000000000", 2841 => "0000000000000000", 2842 => "0000000000000000", 2843 => "0000000000000000", 2844 => "0000000000000000", 2845 => "0000000000000000", 2846 => "0000000000000000", 2847 => "0000000000000000", 2848 => "0000000000000000", 2849 => "0000000000000000", 2850 => "0000000000000000", 2851 => "0000000000000000", 2852 => "0000000000000000", 2853 => "0000000000000000", 2854 => "0000000000000000", 2855 => "0000000000000000", 2856 => "0000000000000000", 2857 => "0000000000000000", 2858 => "0000000000000000", 2859 => "0000000000000000", 2860 => "0000000000000000", 2861 => "0000000000000000", 2862 => "0000000000000000", 2863 => "0000000000000000", 2864 => "0000000000000000", 2865 => "0000000000000000", 2866 => "0000000000000000", 2867 => "0000000000000000", 2868 => "0000000000000000", 2869 => "0000000000000000", 2870 => "0000000000000000", 2871 => "0000000000000000", 2872 => "0000000000000000", 2873 => "0000000000000000", 2874 => "0000000000000000", 2875 => "0000000000000000", 2876 => "0000000000000000", 2877 => "0000000000000000", 2878 => "0000000000000000", 2879 => "0000000000000000", 2880 => "0000000000000000", 2881 => "0000000000000000", 2882 => "0000000000000000", 2883 => "0000000000000000", 2884 => "0000000000000000", 2885 => "0000000000000000", 2886 => "0000000000000000", 2887 => "0000000000000000", 2888 => "0000000000000000", 2889 => "0000000000000000", 2890 => "0000000000000000", 2891 => "0000000000000000", 2892 => "0000000000000000", 2893 => "0000000000000000", 2894 => "0000000000000000", 2895 => "0000000000000000", 2896 => "0000000000000000", 2897 => "0000000000000000", 2898 => "0000000000000000", 2899 => "0000000000000000", 2900 => "0000000000000000", 2901 => "0000000000000000", 2902 => "0000000000000000", 2903 => "0000000000000000", 2904 => "0000000000000000", 2905 => "0000000000000000", 2906 => "0000000000000000", 2907 => "0000000000000000", 2908 => "0000000000000000", 2909 => "0000000000000000", 2910 => "0000000000000000", 2911 => "0000000000000000", 2912 => "0000000000000000", 2913 => "0000000000000000", 2914 => "0000000000000000", 2915 => "0000000000000000", 2916 => "0000000000000000", 2917 => "0000000000000000", 2918 => "0000000000000000", 2919 => "0000000000000000", 2920 => "0000000000000000", 2921 => "0000000000000000", 2922 => "0000000000000000", 2923 => "0000000000000000", 2924 => "0000000000000000", 2925 => "0000000000000000", 2926 => "0000000000000000", 2927 => "0000000000000000", 2928 => "0000000000000000", 2929 => "0000000000000000", 2930 => "0000000000000000", 2931 => "0000000000000000", 2932 => "0000000000000000", 2933 => "0000000000000000", 2934 => "0000000000000000", 2935 => "0000000000000000", 2936 => "0000000000000000", 2937 => "0000000000000000", 2938 => "0000000000000000", 2939 => "0000000000000000", 2940 => "0000000000000000", 2941 => "0000000000000000", 2942 => "0000000000000000", 2943 => "0000000000000000", 2944 => "0000000000000000", 2945 => "0000000000000000", 2946 => "0000000000000000", 2947 => "0000000000000000", 2948 => "0000000000000000", 2949 => "0000000000000000", 2950 => "0000000000000000", 2951 => "0000000000000000", 2952 => "0000000000000000", 2953 => "0000000000000000", 2954 => "0000000000000000", 2955 => "0000000000000000", 2956 => "0000000000000000", 2957 => "0000000000000000", 2958 => "0000000000000000", 2959 => "0000000000000000", 2960 => "0000000000000000", 2961 => "0000000000000000", 2962 => "0000000000000000", 2963 => "0000000000000000", 2964 => "0000000000000000", 2965 => "0000000000000000", 2966 => "0000000000000000", 2967 => "0000000000000000", 2968 => "0000000000000000", 2969 => "0000000000000000", 2970 => "0000000000000000", 2971 => "0000000000000000", 2972 => "0000000000000000", 2973 => "0000000000000000", 2974 => "0000000000000000", 2975 => "0000000000000000", 2976 => "0000000000000000", 2977 => "0000000000000000", 2978 => "0000000000000000", 2979 => "0000000000000000", 2980 => "0000000000000000", 2981 => "0000000000000000", 2982 => "0000000000000000", 2983 => "0000000000000000", 2984 => "0000000000000000", 2985 => "0000000000000000", 2986 => "0000000000000000", 2987 => "0000000000000000", 2988 => "0000000000000000", 2989 => "0000000000000000", 2990 => "0000000000000000", 2991 => "0000000000000000", 2992 => "0000000000000000", 2993 => "0000000000000000", 2994 => "0000000000000000", 2995 => "0000000000000000", 2996 => "0000000000000000", 2997 => "0000000000000000", 2998 => "0000000000000000", 2999 => "0000000000000000", 3000 => "0000000000000000", 3001 => "0000000000000000", 3002 => "0000000000000000", 3003 => "0000000000000000", 3004 => "0000000000000000", 3005 => "0000000000000000", 3006 => "0000000000000000", 3007 => "0000000000000000", 3008 => "0000000000000000", 3009 => "0000000000000000", 3010 => "0000000000000000", 3011 => "0000000000000000", 3012 => "0000000000000000", 3013 => "0000000000000000", 3014 => "0000000000000000", 3015 => "0000000000000000", 3016 => "0000000000000000", 3017 => "0000000000000000", 3018 => "0000000000000000", 3019 => "0000000000000000", 3020 => "0000000000000000", 3021 => "0000000000000000", 3022 => "0000000000000000", 3023 => "0000000000000000", 3024 => "0000000000000000", 3025 => "0000000000000000", 3026 => "0000000000000000", 3027 => "0000000000000000", 3028 => "0000000000000000", 3029 => "0000000000000000", 3030 => "0000000000000000", 3031 => "0000000000000000", 3032 => "0000000000000000", 3033 => "0000000000000000", 3034 => "0000000000000000", 3035 => "0000000000000000", 3036 => "0000000000000000", 3037 => "0000000000000000", 3038 => "0000000000000000", 3039 => "0000000000000000", 3040 => "0000000000000000", 3041 => "0000000000000000", 3042 => "0000000000000000", 3043 => "0000000000000000", 3044 => "0000000000000000", 3045 => "0000000000000000", 3046 => "0000000000000000", 3047 => "0000000000000000", 3048 => "0000000000000000", 3049 => "0000000000000000", 3050 => "0000000000000000", 3051 => "0000000000000000", 3052 => "0000000000000000", 3053 => "0000000000000000", 3054 => "0000000000000000", 3055 => "0000000000000000", 3056 => "0000000000000000", 3057 => "0000000000000000", 3058 => "0000000000000000", 3059 => "0000000000000000", 3060 => "0000000000000000", 3061 => "0000000000000000", 3062 => "0000000000000000", 3063 => "0000000000000000", 3064 => "0000000000000000", 3065 => "0000000000000000", 3066 => "0000000000000000", 3067 => "0000000000000000", 3068 => "0000000000000000", 3069 => "0000000000000000", 3070 => "0000000000000000", 3071 => "0000000000000000", 3072 => "0000000000000000", 3073 => "0000000000000000", 3074 => "0000000000000000", 3075 => "0000000000000000", 3076 => "0000000000000000", 3077 => "0000000000000000", 3078 => "0000000000000000", 3079 => "0000000000000000", 3080 => "0000000000000000", 3081 => "0000000000000000", 3082 => "0000000000000000", 3083 => "0000000000000000", 3084 => "0000000000000000", 3085 => "0000000000000000", 3086 => "0000000000000000", 3087 => "0000000000000000", 3088 => "0000000000000000", 3089 => "0000000000000000", 3090 => "0000000000000000", 3091 => "0000000000000000", 3092 => "0000000000000000", 3093 => "0000000000000000", 3094 => "0000000000000000", 3095 => "0000000000000000", 3096 => "0000000000000000", 3097 => "0000000000000000", 3098 => "0000000000000000", 3099 => "0000000000000000", 3100 => "0000000000000000", 3101 => "0000000000000000", 3102 => "0000000000000000", 3103 => "0000000000000000", 3104 => "0000000000000000", 3105 => "0000000000000000", 3106 => "0000000000000000", 3107 => "0000000000000000", 3108 => "0000000000000000", 3109 => "0000000000000000", 3110 => "0000000000000000", 3111 => "0000000000000000", 3112 => "0000000000000000", 3113 => "0000000000000000", 3114 => "0000000000000000", 3115 => "0000000000000000", 3116 => "0000000000000000", 3117 => "0000000000000000", 3118 => "0000000000000000", 3119 => "0000000000000000", 3120 => "0000000000000000", 3121 => "0000000000000000", 3122 => "0000000000000000", 3123 => "0000000000000000", 3124 => "0000000000000000", 3125 => "0000000000000000", 3126 => "0000000000000000", 3127 => "0000000000000000", 3128 => "0000000000000000", 3129 => "0000000000000000", 3130 => "0000000000000000", 3131 => "0000000000000000", 3132 => "0000000000000000", 3133 => "0000000000000000", 3134 => "0000000000000000", 3135 => "0000000000000000", 3136 => "0000000000000000", 3137 => "0000000000000000", 3138 => "0000000000000000", 3139 => "0000000000000000", 3140 => "0000000000000000", 3141 => "0000000000000000", 3142 => "0000000000000000", 3143 => "0000000000000000", 3144 => "0000000000000000", 3145 => "0000000000000000", 3146 => "0000000000000000", 3147 => "0000000000000000", 3148 => "0000000000000000", 3149 => "0000000000000000", 3150 => "0000000000000000", 3151 => "0000000000000000", 3152 => "0000000000000000", 3153 => "0000000000000000", 3154 => "0000000000000000", 3155 => "0000000000000000", 3156 => "0000000000000000", 3157 => "0000000000000000", 3158 => "0000000000000000", 3159 => "0000000000000000", 3160 => "0000000000000000", 3161 => "0000000000000000", 3162 => "0000000000000000", 3163 => "0000000000000000", 3164 => "0000000000000000", 3165 => "0000000000000000", 3166 => "0000000000000000", 3167 => "0000000000000000", 3168 => "0000000000000000", 3169 => "0000000000000000", 3170 => "0000000000000000", 3171 => "0000000000000000", 3172 => "0000000000000000", 3173 => "0000000000000000", 3174 => "0000000000000000", 3175 => "0000000000000000", 3176 => "0000000000000000", 3177 => "0000000000000000", 3178 => "0000000000000000", 3179 => "0000000000000000", 3180 => "0000000000000000", 3181 => "0000000000000000", 3182 => "0000000000000000", 3183 => "0000000000000000", 3184 => "0000000000000000", 3185 => "0000000000000000", 3186 => "0000000000000000", 3187 => "0000000000000000", 3188 => "0000000000000000", 3189 => "0000000000000000", 3190 => "0000000000000000", 3191 => "0000000000000000", 3192 => "0000000000000000", 3193 => "0000000000000000", 3194 => "0000000000000000", 3195 => "0000000000000000", 3196 => "0000000000000000", 3197 => "0000000000000000", 3198 => "0000000000000000", 3199 => "0000000000000000", 3200 => "0000000000000000", 3201 => "0000000000000000", 3202 => "0000000000000000", 3203 => "0000000000000000", 3204 => "0000000000000000", 3205 => "0000000000000000", 3206 => "0000000000000000", 3207 => "0000000000000000", 3208 => "0000000000000000", 3209 => "0000000000000000", 3210 => "0000000000000000", 3211 => "0000000000000000", 3212 => "0000000000000000", 3213 => "0000000000000000", 3214 => "0000000000000000", 3215 => "0000000000000000", 3216 => "0000000000000000", 3217 => "0000000000000000", 3218 => "0000000000000000", 3219 => "0000000000000000", 3220 => "0000000000000000", 3221 => "0000000000000000", 3222 => "0000000000000000", 3223 => "0000000000000000", 3224 => "0000000000000000", 3225 => "0000000000000000", 3226 => "0000000000000000", 3227 => "0000000000000000", 3228 => "0000000000000000", 3229 => "0000000000000000", 3230 => "0000000000000000", 3231 => "0000000000000000", 3232 => "0000000000000000", 3233 => "0000000000000000", 3234 => "0000000000000000", 3235 => "0000000000000000", 3236 => "0000000000000000", 3237 => "0000000000000000", 3238 => "0000000000000000", 3239 => "0000000000000000", 3240 => "0000000000000000", 3241 => "0000000000000000", 3242 => "0000000000000000", 3243 => "0000000000000000", 3244 => "0000000000000000", 3245 => "0000000000000000", 3246 => "0000000000000000", 3247 => "0000000000000000", 3248 => "0000000000000000", 3249 => "0000000000000000", 3250 => "0000000000000000", 3251 => "0000000000000000", 3252 => "0000000000000000", 3253 => "0000000000000000", 3254 => "0000000000000000", 3255 => "0000000000000000", 3256 => "0000000000000000", 3257 => "0000000000000000", 3258 => "0000000000000000", 3259 => "0000000000000000", 3260 => "0000000000000000", 3261 => "0000000000000000", 3262 => "0000000000000000", 3263 => "0000000000000000", 3264 => "0000000000000000", 3265 => "0000000000000000", 3266 => "0000000000000000", 3267 => "0000000000000000", 3268 => "0000000000000000", 3269 => "0000000000000000", 3270 => "0000000000000000", 3271 => "0000000000000000", 3272 => "0000000000000000", 3273 => "0000000000000000", 3274 => "0000000000000000", 3275 => "0000000000000000", 3276 => "0000000000000000", 3277 => "0000000000000000", 3278 => "0000000000000000", 3279 => "0000000000000000", 3280 => "0000000000000000", 3281 => "0000000000000000", 3282 => "0000000000000000", 3283 => "0000000000000000", 3284 => "0000000000000000", 3285 => "0000000000000000", 3286 => "0000000000000000", 3287 => "0000000000000000", 3288 => "0000000000000000", 3289 => "0000000000000000", 3290 => "0000000000000000", 3291 => "0000000000000000", 3292 => "0000000000000000", 3293 => "0000000000000000", 3294 => "0000000000000000", 3295 => "0000000000000000", 3296 => "0000000000000000", 3297 => "0000000000000000", 3298 => "0000000000000000", 3299 => "0000000000000000", 3300 => "0000000000000000", 3301 => "0000000000000000", 3302 => "0000000000000000", 3303 => "0000000000000000", 3304 => "0000000000000000", 3305 => "0000000000000000", 3306 => "0000000000000000", 3307 => "0000000000000000", 3308 => "0000000000000000", 3309 => "0000000000000000", 3310 => "0000000000000000", 3311 => "0000000000000000", 3312 => "0000000000000000", 3313 => "0000000000000000", 3314 => "0000000000000000", 3315 => "0000000000000000", 3316 => "0000000000000000", 3317 => "0000000000000000", 3318 => "0000000000000000", 3319 => "0000000000000000", 3320 => "0000000000000000", 3321 => "0000000000000000", 3322 => "0000000000000000", 3323 => "0000000000000000", 3324 => "0000000000000000", 3325 => "0000000000000000", 3326 => "0000000000000000", 3327 => "0000000000000000", 3328 => "0000000000000000", 3329 => "0000000000000000", 3330 => "0000000000000000", 3331 => "0000000000000000", 3332 => "0000000000000000", 3333 => "0000000000000000", 3334 => "0000000000000000", 3335 => "0000000000000000", 3336 => "0000000000000000", 3337 => "0000000000000000", 3338 => "0000000000000000", 3339 => "0000000000000000", 3340 => "0000000000000000", 3341 => "0000000000000000", 3342 => "0000000000000000", 3343 => "0000000000000000", 3344 => "0000000000000000", 3345 => "0000000000000000", 3346 => "0000000000000000", 3347 => "0000000000000000", 3348 => "0000000000000000", 3349 => "0000000000000000", 3350 => "0000000000000000", 3351 => "0000000000000000", 3352 => "0000000000000000", 3353 => "0000000000000000", 3354 => "0000000000000000", 3355 => "0000000000000000", 3356 => "0000000000000000", 3357 => "0000000000000000", 3358 => "0000000000000000", 3359 => "0000000000000000", 3360 => "0000000000000000", 3361 => "0000000000000000", 3362 => "0000000000000000", 3363 => "0000000000000000", 3364 => "0000000000000000", 3365 => "0000000000000000", 3366 => "0000000000000000", 3367 => "0000000000000000", 3368 => "0000000000000000", 3369 => "0000000000000000", 3370 => "0000000000000000", 3371 => "0000000000000000", 3372 => "0000000000000000", 3373 => "0000000000000000", 3374 => "0000000000000000", 3375 => "0000000000000000", 3376 => "0000000000000000", 3377 => "0000000000000000", 3378 => "0000000000000000", 3379 => "0000000000000000", 3380 => "0000000000000000", 3381 => "0000000000000000", 3382 => "0000000000000000", 3383 => "0000000000000000", 3384 => "0000000000000000", 3385 => "0000000000000000", 3386 => "0000000000000000", 3387 => "0000000000000000", 3388 => "0000000000000000", 3389 => "0000000000000000", 3390 => "0000000000000000", 3391 => "0000000000000000", 3392 => "0000000000000000", 3393 => "0000000000000000", 3394 => "0000000000000000", 3395 => "0000000000000000", 3396 => "0000000000000000", 3397 => "0000000000000000", 3398 => "0000000000000000", 3399 => "0000000000000000", 3400 => "0000000000000000", 3401 => "0000000000000000", 3402 => "0000000000000000", 3403 => "0000000000000000", 3404 => "0000000000000000", 3405 => "0000000000000000", 3406 => "0000000000000000", 3407 => "0000000000000000", 3408 => "0000000000000000", 3409 => "0000000000000000", 3410 => "0000000000000000", 3411 => "0000000000000000", 3412 => "0000000000000000", 3413 => "0000000000000000", 3414 => "0000000000000000", 3415 => "0000000000000000", 3416 => "0000000000000000", 3417 => "0000000000000000", 3418 => "0000000000000000", 3419 => "0000000000000000", 3420 => "0000000000000000", 3421 => "0000000000000000", 3422 => "0000000000000000", 3423 => "0000000000000000", 3424 => "0000000000000000", 3425 => "0000000000000000", 3426 => "0000000000000000", 3427 => "0000000000000000", 3428 => "0000000000000000", 3429 => "0000000000000000", 3430 => "0000000000000000", 3431 => "0000000000000000", 3432 => "0000000000000000", 3433 => "0000000000000000", 3434 => "0000000000000000", 3435 => "0000000000000000", 3436 => "0000000000000000", 3437 => "0000000000000000", 3438 => "0000000000000000", 3439 => "0000000000000000", 3440 => "0000000000000000", 3441 => "0000000000000000", 3442 => "0000000000000000", 3443 => "0000000000000000", 3444 => "0000000000000000", 3445 => "0000000000000000", 3446 => "0000000000000000", 3447 => "0000000000000000", 3448 => "0000000000000000", 3449 => "0000000000000000", 3450 => "0000000000000000", 3451 => "0000000000000000", 3452 => "0000000000000000", 3453 => "0000000000000000", 3454 => "0000000000000000", 3455 => "0000000000000000", 3456 => "0000000000000000", 3457 => "0000000000000000", 3458 => "0000000000000000", 3459 => "0000000000000000", 3460 => "0000000000000000", 3461 => "0000000000000000", 3462 => "0000000000000000", 3463 => "0000000000000000", 3464 => "0000000000000000", 3465 => "0000000000000000", 3466 => "0000000000000000", 3467 => "0000000000000000", 3468 => "0000000000000000", 3469 => "0000000000000000", 3470 => "0000000000000000", 3471 => "0000000000000000", 3472 => "0000000000000000", 3473 => "0000000000000000", 3474 => "0000000000000000", 3475 => "0000000000000000", 3476 => "0000000000000000", 3477 => "0000000000000000", 3478 => "0000000000000000", 3479 => "0000000000000000", 3480 => "0000000000000000", 3481 => "0000000000000000", 3482 => "0000000000000000", 3483 => "0000000000000000", 3484 => "0000000000000000", 3485 => "0000000000000000", 3486 => "0000000000000000", 3487 => "0000000000000000", 3488 => "0000000000000000", 3489 => "0000000000000000", 3490 => "0000000000000000", 3491 => "0000000000000000", 3492 => "0000000000000000", 3493 => "0000000000000000", 3494 => "0000000000000000", 3495 => "0000000000000000", 3496 => "0000000000000000", 3497 => "0000000000000000", 3498 => "0000000000000000", 3499 => "0000000000000000", 3500 => "0000000000000000", 3501 => "0000000000000000", 3502 => "0000000000000000", 3503 => "0000000000000000", 3504 => "0000000000000000", 3505 => "0000000000000000", 3506 => "0000000000000000", 3507 => "0000000000000000", 3508 => "0000000000000000", 3509 => "0000000000000000", 3510 => "0000000000000000", 3511 => "0000000000000000", 3512 => "0000000000000000", 3513 => "0000000000000000", 3514 => "0000000000000000", 3515 => "0000000000000000", 3516 => "0000000000000000", 3517 => "0000000000000000", 3518 => "0000000000000000", 3519 => "0000000000000000", 3520 => "0000000000000000", 3521 => "0000000000000000", 3522 => "0000000000000000", 3523 => "0000000000000000", 3524 => "0000000000000000", 3525 => "0000000000000000", 3526 => "0000000000000000", 3527 => "0000000000000000", 3528 => "0000000000000000", 3529 => "0000000000000000", 3530 => "0000000000000000", 3531 => "0000000000000000", 3532 => "0000000000000000", 3533 => "0000000000000000", 3534 => "0000000000000000", 3535 => "0000000000000000", 3536 => "0000000000000000", 3537 => "0000000000000000", 3538 => "0000000000000000", 3539 => "0000000000000000", 3540 => "0000000000000000", 3541 => "0000000000000000", 3542 => "0000000000000000", 3543 => "0000000000000000", 3544 => "0000000000000000", 3545 => "0000000000000000", 3546 => "0000000000000000", 3547 => "0000000000000000", 3548 => "0000000000000000", 3549 => "0000000000000000", 3550 => "0000000000000000", 3551 => "0000000000000000", 3552 => "0000000000000000", 3553 => "0000000000000000", 3554 => "0000000000000000", 3555 => "0000000000000000", 3556 => "0000000000000000", 3557 => "0000000000000000", 3558 => "0000000000000000", 3559 => "0000000000000000", 3560 => "0000000000000000", 3561 => "0000000000000000", 3562 => "0000000000000000", 3563 => "0000000000000000", 3564 => "0000000000000000", 3565 => "0000000000000000", 3566 => "0000000000000000", 3567 => "0000000000000000", 3568 => "0000000000000000", 3569 => "0000000000000000", 3570 => "0000000000000000", 3571 => "0000000000000000", 3572 => "0000000000000000", 3573 => "0000000000000000", 3574 => "0000000000000000", 3575 => "0000000000000000", 3576 => "0000000000000000", 3577 => "0000000000000000", 3578 => "0000000000000000", 3579 => "0000000000000000", 3580 => "0000000000000000", 3581 => "0000000000000000", 3582 => "0000000000000000", 3583 => "0000000000000000", 3584 => "0000000000000000", 3585 => "0000000000000000", 3586 => "0000000000000000", 3587 => "0000000000000000", 3588 => "0000000000000000", 3589 => "0000000000000000", 3590 => "0000000000000000", 3591 => "0000000000000000", 3592 => "0000000000000000", 3593 => "0000000000000000", 3594 => "0000000000000000", 3595 => "0000000000000000", 3596 => "0000000000000000", 3597 => "0000000000000000", 3598 => "0000000000000000", 3599 => "0000000000000000", 3600 => "0000000000000000", 3601 => "0000000000000000", 3602 => "0000000000000000", 3603 => "0000000000000000", 3604 => "0000000000000000", 3605 => "0000000000000000", 3606 => "0000000000000000", 3607 => "0000000000000000", 3608 => "0000000000000000", 3609 => "0000000000000000", 3610 => "0000000000000000", 3611 => "0000000000000000", 3612 => "0000000000000000", 3613 => "0000000000000000", 3614 => "0000000000000000", 3615 => "0000000000000000", 3616 => "0000000000000000", 3617 => "0000000000000000", 3618 => "0000000000000000", 3619 => "0000000000000000", 3620 => "0000000000000000", 3621 => "0000000000000000", 3622 => "0000000000000000", 3623 => "0000000000000000", 3624 => "0000000000000000", 3625 => "0000000000000000", 3626 => "0000000000000000", 3627 => "0000000000000000", 3628 => "0000000000000000", 3629 => "0000000000000000", 3630 => "0000000000000000", 3631 => "0000000000000000", 3632 => "0000000000000000", 3633 => "0000000000000000", 3634 => "0000000000000000", 3635 => "0000000000000000", 3636 => "0000000000000000", 3637 => "0000000000000000", 3638 => "0000000000000000", 3639 => "0000000000000000", 3640 => "0000000000000000", 3641 => "0000000000000000", 3642 => "0000000000000000", 3643 => "0000000000000000", 3644 => "0000000000000000", 3645 => "0000000000000000", 3646 => "0000000000000000", 3647 => "0000000000000000", 3648 => "0000000000000000", 3649 => "0000000000000000", 3650 => "0000000000000000", 3651 => "0000000000000000", 3652 => "0000000000000000", 3653 => "0000000000000000", 3654 => "0000000000000000", 3655 => "0000000000000000", 3656 => "0000000000000000", 3657 => "0000000000000000", 3658 => "0000000000000000", 3659 => "0000000000000000", 3660 => "0000000000000000", 3661 => "0000000000000000", 3662 => "0000000000000000", 3663 => "0000000000000000", 3664 => "0000000000000000", 3665 => "0000000000000000", 3666 => "0000000000000000", 3667 => "0000000000000000", 3668 => "0000000000000000", 3669 => "0000000000000000", 3670 => "0000000000000000", 3671 => "0000000000000000", 3672 => "0000000000000000", 3673 => "0000000000000000", 3674 => "0000000000000000", 3675 => "0000000000000000", 3676 => "0000000000000000", 3677 => "0000000000000000", 3678 => "0000000000000000", 3679 => "0000000000000000", 3680 => "0000000000000000", 3681 => "0000000000000000", 3682 => "0000000000000000", 3683 => "0000000000000000", 3684 => "0000000000000000", 3685 => "0000000000000000", 3686 => "0000000000000000", 3687 => "0000000000000000", 3688 => "0000000000000000", 3689 => "0000000000000000", 3690 => "0000000000000000", 3691 => "0000000000000000", 3692 => "0000000000000000", 3693 => "0000000000000000", 3694 => "0000000000000000", 3695 => "0000000000000000", 3696 => "0000000000000000", 3697 => "0000000000000000", 3698 => "0000000000000000", 3699 => "0000000000000000", 3700 => "0000000000000000", 3701 => "0000000000000000", 3702 => "0000000000000000", 3703 => "0000000000000000", 3704 => "0000000000000000", 3705 => "0000000000000000", 3706 => "0000000000000000", 3707 => "0000000000000000", 3708 => "0000000000000000", 3709 => "0000000000000000", 3710 => "0000000000000000", 3711 => "0000000000000000", 3712 => "0000000000000000", 3713 => "0000000000000000", 3714 => "0000000000000000", 3715 => "0000000000000000", 3716 => "0000000000000000", 3717 => "0000000000000000", 3718 => "0000000000000000", 3719 => "0000000000000000", 3720 => "0000000000000000", 3721 => "0000000000000000", 3722 => "0000000000000000", 3723 => "0000000000000000", 3724 => "0000000000000000", 3725 => "0000000000000000", 3726 => "0000000000000000", 3727 => "0000000000000000", 3728 => "0000000000000000", 3729 => "0000000000000000", 3730 => "0000000000000000", 3731 => "0000000000000000", 3732 => "0000000000000000", 3733 => "0000000000000000", 3734 => "0000000000000000", 3735 => "0000000000000000", 3736 => "0000000000000000", 3737 => "0000000000000000", 3738 => "0000000000000000", 3739 => "0000000000000000", 3740 => "0000000000000000", 3741 => "0000000000000000", 3742 => "0000000000000000", 3743 => "0000000000000000", 3744 => "0000000000000000", 3745 => "0000000000000000", 3746 => "0000000000000000", 3747 => "0000000000000000", 3748 => "0000000000000000", 3749 => "0000000000000000", 3750 => "0000000000000000", 3751 => "0000000000000000", 3752 => "0000000000000000", 3753 => "0000000000000000", 3754 => "0000000000000000", 3755 => "0000000000000000", 3756 => "0000000000000000", 3757 => "0000000000000000", 3758 => "0000000000000000", 3759 => "0000000000000000", 3760 => "0000000000000000", 3761 => "0000000000000000", 3762 => "0000000000000000", 3763 => "0000000000000000", 3764 => "0000000000000000", 3765 => "0000000000000000", 3766 => "0000000000000000", 3767 => "0000000000000000", 3768 => "0000000000000000", 3769 => "0000000000000000", 3770 => "0000000000000000", 3771 => "0000000000000000", 3772 => "0000000000000000", 3773 => "0000000000000000", 3774 => "0000000000000000", 3775 => "0000000000000000", 3776 => "0000000000000000", 3777 => "0000000000000000", 3778 => "0000000000000000", 3779 => "0000000000000000", 3780 => "0000000000000000", 3781 => "0000000000000000", 3782 => "0000000000000000", 3783 => "0000000000000000", 3784 => "0000000000000000", 3785 => "0000000000000000", 3786 => "0000000000000000", 3787 => "0000000000000000", 3788 => "0000000000000000", 3789 => "0000000000000000", 3790 => "0000000000000000", 3791 => "0000000000000000", 3792 => "0000000000000000", 3793 => "0000000000000000", 3794 => "0000000000000000", 3795 => "0000000000000000", 3796 => "0000000000000000", 3797 => "0000000000000000", 3798 => "0000000000000000", 3799 => "0000000000000000", 3800 => "0000000000000000", 3801 => "0000000000000000", 3802 => "0000000000000000", 3803 => "0000000000000000", 3804 => "0000000000000000", 3805 => "0000000000000000", 3806 => "0000000000000000", 3807 => "0000000000000000", 3808 => "0000000000000000", 3809 => "0000000000000000", 3810 => "0000000000000000", 3811 => "0000000000000000", 3812 => "0000000000000000", 3813 => "0000000000000000", 3814 => "0000000000000000", 3815 => "0000000000000000", 3816 => "0000000000000000", 3817 => "0000000000000000", 3818 => "0000000000000000", 3819 => "0000000000000000", 3820 => "0000000000000000", 3821 => "0000000000000000", 3822 => "0000000000000000", 3823 => "0000000000000000", 3824 => "0000000000000000", 3825 => "0000000000000000", 3826 => "0000000000000000", 3827 => "0000000000000000", 3828 => "0000000000000000", 3829 => "0000000000000000", 3830 => "0000000000000000", 3831 => "0000000000000000", 3832 => "0000000000000000", 3833 => "0000000000000000", 3834 => "0000000000000000", 3835 => "0000000000000000", 3836 => "0000000000000000", 3837 => "0000000000000000", 3838 => "0000000000000000", 3839 => "0000000000000000", 3840 => "0000000000000000", 3841 => "0000000000000000", 3842 => "0000000000000000", 3843 => "0000000000000000", 3844 => "0000000000000000", 3845 => "0000000000000000", 3846 => "0000000000000000", 3847 => "0000000000000000", 3848 => "0000000000000000", 3849 => "0000000000000000", 3850 => "0000000000000000", 3851 => "0000000000000000", 3852 => "0000000000000000", 3853 => "0000000000000000", 3854 => "0000000000000000", 3855 => "0000000000000000", 3856 => "0000000000000000", 3857 => "0000000000000000", 3858 => "0000000000000000", 3859 => "0000000000000000", 3860 => "0000000000000000", 3861 => "0000000000000000", 3862 => "0000000000000000", 3863 => "0000000000000000", 3864 => "0000000000000000", 3865 => "0000000000000000", 3866 => "0000000000000000", 3867 => "0000000000000000", 3868 => "0000000000000000", 3869 => "0000000000000000", 3870 => "0000000000000000", 3871 => "0000000000000000", 3872 => "0000000000000000", 3873 => "0000000000000000", 3874 => "0000000000000000", 3875 => "0000000000000000", 3876 => "0000000000000000", 3877 => "0000000000000000", 3878 => "0000000000000000", 3879 => "0000000000000000", 3880 => "0000000000000000", 3881 => "0000000000000000", 3882 => "0000000000000000", 3883 => "0000000000000000", 3884 => "0000000000000000", 3885 => "0000000000000000", 3886 => "0000000000000000", 3887 => "0000000000000000", 3888 => "0000000000000000", 3889 => "0000000000000000", 3890 => "0000000000000000", 3891 => "0000000000000000", 3892 => "0000000000000000", 3893 => "0000000000000000", 3894 => "0000000000000000", 3895 => "0000000000000000", 3896 => "0000000000000000", 3897 => "0000000000000000", 3898 => "0000000000000000", 3899 => "0000000000000000", 3900 => "0000000000000000", 3901 => "0000000000000000", 3902 => "0000000000000000", 3903 => "0000000000000000", 3904 => "0000000000000000", 3905 => "0000000000000000", 3906 => "0000000000000000", 3907 => "0000000000000000", 3908 => "0000000000000000", 3909 => "0000000000000000", 3910 => "0000000000000000", 3911 => "0000000000000000", 3912 => "0000000000000000", 3913 => "0000000000000000", 3914 => "0000000000000000", 3915 => "0000000000000000", 3916 => "0000000000000000", 3917 => "0000000000000000", 3918 => "0000000000000000", 3919 => "0000000000000000", 3920 => "0000000000000000", 3921 => "0000000000000000", 3922 => "0000000000000000", 3923 => "0000000000000000", 3924 => "0000000000000000", 3925 => "0000000000000000", 3926 => "0000000000000000", 3927 => "0000000000000000", 3928 => "0000000000000000", 3929 => "0000000000000000", 3930 => "0000000000000000", 3931 => "0000000000000000", 3932 => "0000000000000000", 3933 => "0000000000000000", 3934 => "0000000000000000", 3935 => "0000000000000000", 3936 => "0000000000000000", 3937 => "0000000000000000", 3938 => "0000000000000000", 3939 => "0000000000000000", 3940 => "0000000000000000", 3941 => "0000000000000000", 3942 => "0000000000000000", 3943 => "0000000000000000", 3944 => "0000000000000000", 3945 => "0000000000000000", 3946 => "0000000000000000", 3947 => "0000000000000000", 3948 => "0000000000000000", 3949 => "0000000000000000", 3950 => "0000000000000000", 3951 => "0000000000000000", 3952 => "0000000000000000", 3953 => "0000000000000000", 3954 => "0000000000000000", 3955 => "0000000000000000", 3956 => "0000000000000000", 3957 => "0000000000000000", 3958 => "0000000000000000", 3959 => "0000000000000000", 3960 => "0000000000000000", 3961 => "0000000000000000", 3962 => "0000000000000000", 3963 => "0000000000000000", 3964 => "0000000000000000", 3965 => "0000000000000000", 3966 => "0000000000000000", 3967 => "0000000000000000", 3968 => "0000000000000000", 3969 => "0000000000000000", 3970 => "0000000000000000", 3971 => "0000000000000000", 3972 => "0000000000000000", 3973 => "0000000000000000", 3974 => "0000000000000000", 3975 => "0000000000000000", 3976 => "0000000000000000", 3977 => "0000000000000000", 3978 => "0000000000000000", 3979 => "0000000000000000", 3980 => "0000000000000000", 3981 => "0000000000000000", 3982 => "0000000000000000", 3983 => "0000000000000000", 3984 => "0000000000000000", 3985 => "0000000000000000", 3986 => "0000000000000000", 3987 => "0000000000000000", 3988 => "0000000000000000", 3989 => "0000000000000000", 3990 => "0000000000000000", 3991 => "0000000000000000", 3992 => "0000000000000000", 3993 => "0000000000000000", 3994 => "0000000000000000", 3995 => "0000000000000000", 3996 => "0000000000000000", 3997 => "0000000000000000", 3998 => "0000000000000000", 3999 => "0000000000000000", 4000 => "0000000000000000", 4001 => "0000000000000000", 4002 => "0000000000000000", 4003 => "0000000000000000", 4004 => "0000000000000000", 4005 => "0000000000000000", 4006 => "0000000000000000", 4007 => "0000000000000000", 4008 => "0000000000000000", 4009 => "0000000000000000", 4010 => "0000000000000000", 4011 => "0000000000000000", 4012 => "0000000000000000", 4013 => "0000000000000000", 4014 => "0000000000000000", 4015 => "0000000000000000", 4016 => "0000000000000000", 4017 => "0000000000000000", 4018 => "0000000000000000", 4019 => "0000000000000000", 4020 => "0000000000000000", 4021 => "0000000000000000", 4022 => "0000000000000000", 4023 => "0000000000000000", 4024 => "0000000000000000", 4025 => "0000000000000000", 4026 => "0000000000000000", 4027 => "0000000000000000", 4028 => "0000000000000000", 4029 => "0000000000000000", 4030 => "0000000000000000", 4031 => "0000000000000000", 4032 => "0000000000000000", 4033 => "0000000000000000", 4034 => "0000000000000000", 4035 => "0000000000000000", 4036 => "0000000000000000", 4037 => "0000000000000000", 4038 => "0000000000000000", 4039 => "0000000000000000", 4040 => "0000000000000000", 4041 => "0000000000000000", 4042 => "0000000000000000", 4043 => "0000000000000000", 4044 => "0000000000000000", 4045 => "0000000000000000", 4046 => "0000000000000000", 4047 => "0000000000000000", 4048 => "0000000000000000", 4049 => "0000000000000000", 4050 => "0000000000000000", 4051 => "0000000000000000", 4052 => "0000000000000000", 4053 => "0000000000000000", 4054 => "0000000000000000", 4055 => "0000000000000000", 4056 => "0000000000000000", 4057 => "0000000000000000", 4058 => "0000000000000000", 4059 => "0000000000000000", 4060 => "0000000000000000", 4061 => "0000000000000000", 4062 => "0000000000000000", 4063 => "0000000000000000", 4064 => "0000000000000000", 4065 => "0000000000000000", 4066 => "0000000000000000", 4067 => "0000000000000000", 4068 => "0000000000000000", 4069 => "0000000000000000", 4070 => "0000000000000000", 4071 => "0000000000000000", 4072 => "0000000000000000", 4073 => "0000000000000000", 4074 => "0000000000000000", 4075 => "0000000000000000", 4076 => "0000000000000000", 4077 => "0000000000000000", 4078 => "0000000000000000", 4079 => "0000000000000000", 4080 => "0000000000000000", 4081 => "0000000000000000", 4082 => "0000000000000000", 4083 => "0000000000000000", 4084 => "0000000000000000", 4085 => "0000000000000000", 4086 => "0000000000000000", 4087 => "0000000000000000", 4088 => "0000000000000000", 4089 => "0000000000000000", 4090 => "0000000000000000", 4091 => "0000000000000000", 4092 => "0000000000000000", 4093 => "0000000000000000", 4094 => "0000000000000000", 4095 => "0000000000000000", 4096 => "0000000000000000", 4097 => "0000000000000000", 4098 => "0000000000000000", 4099 => "0000000000000000", 4100 => "0000000000000000", 4101 => "0000000000000000", 4102 => "0000000000000000", 4103 => "0000000000000000", 4104 => "0000000000000000", 4105 => "0000000000000000", 4106 => "0000000000000000", 4107 => "0000000000000000", 4108 => "0000000000000000", 4109 => "0000000000000000", 4110 => "0000000000000000", 4111 => "0000000000000000", 4112 => "0000000000000000", 4113 => "0000000000000000", 4114 => "0000000000000000", 4115 => "0000000000000000", 4116 => "0000000000000000", 4117 => "0000000000000000", 4118 => "0000000000000000", 4119 => "0000000000000000", 4120 => "0000000000000000", 4121 => "0000000000000000", 4122 => "0000000000000000", 4123 => "0000000000000000", 4124 => "0000000000000000", 4125 => "0000000000000000", 4126 => "0000000000000000", 4127 => "0000000000000000", 4128 => "0000000000000000", 4129 => "0000000000000000", 4130 => "0000000000000000", 4131 => "0000000000000000", 4132 => "0000000000000000", 4133 => "0000000000000000", 4134 => "0000000000000000", 4135 => "0000000000000000", 4136 => "0000000000000000", 4137 => "0000000000000000", 4138 => "0000000000000000", 4139 => "0000000000000000", 4140 => "0000000000000000", 4141 => "0000000000000000", 4142 => "0000000000000000", 4143 => "0000000000000000", 4144 => "0000000000000000", 4145 => "0000000000000000", 4146 => "0000000000000000", 4147 => "0000000000000000", 4148 => "0000000000000000", 4149 => "0000000000000000", 4150 => "0000000000000000", 4151 => "0000000000000000", 4152 => "0000000000000000", 4153 => "0000000000000000", 4154 => "0000000000000000", 4155 => "0000000000000000", 4156 => "0000000000000000", 4157 => "0000000000000000", 4158 => "0000000000000000", 4159 => "0000000000000000", 4160 => "0000000000000000", 4161 => "0000000000000000", 4162 => "0000000000000000", 4163 => "0000000000000000", 4164 => "0000000000000000", 4165 => "0000000000000000", 4166 => "0000000000000000", 4167 => "0000000000000000", 4168 => "0000000000000000", 4169 => "0000000000000000", 4170 => "0000000000000000", 4171 => "0000000000000000", 4172 => "0000000000000000", 4173 => "0000000000000000", 4174 => "0000000000000000", 4175 => "0000000000000000", 4176 => "0000000000000000", 4177 => "0000000000000000", 4178 => "0000000000000000", 4179 => "0000000000000000", 4180 => "0000000000000000", 4181 => "0000000000000000", 4182 => "0000000000000000", 4183 => "0000000000000000", 4184 => "0000000000000000", 4185 => "0000000000000000", 4186 => "0000000000000000", 4187 => "0000000000000000", 4188 => "0000000000000000", 4189 => "0000000000000000", 4190 => "0000000000000000", 4191 => "0000000000000000", 4192 => "0000000000000000", 4193 => "0000000000000000", 4194 => "0000000000000000", 4195 => "0000000000000000", 4196 => "0000000000000000", 4197 => "0000000000000000", 4198 => "0000000000000000", 4199 => "0000000000000000", 4200 => "0000000000000000", 4201 => "0000000000000000", 4202 => "0000000000000000", 4203 => "0000000000000000", 4204 => "0000000000000000", 4205 => "0000000000000000", 4206 => "0000000000000000", 4207 => "0000000000000000", 4208 => "0000000000000000", 4209 => "0000000000000000", 4210 => "0000000000000000", 4211 => "0000000000000000", 4212 => "0000000000000000", 4213 => "0000000000000000", 4214 => "0000000000000000", 4215 => "0000000000000000", 4216 => "0000000000000000", 4217 => "0000000000000000", 4218 => "0000000000000000", 4219 => "0000000000000000", 4220 => "0000000000000000", 4221 => "0000000000000000", 4222 => "0000000000000000", 4223 => "0000000000000000", 4224 => "0000000000000000", 4225 => "0000000000000000", 4226 => "0000000000000000", 4227 => "0000000000000000", 4228 => "0000000000000000", 4229 => "0000000000000000", 4230 => "0000000000000000", 4231 => "0000000000000000", 4232 => "0000000000000000", 4233 => "0000000000000000", 4234 => "0000000000000000", 4235 => "0000000000000000", 4236 => "0000000000000000", 4237 => "0000000000000000", 4238 => "0000000000000000", 4239 => "0000000000000000", 4240 => "0000000000000000", 4241 => "0000000000000000", 4242 => "0000000000000000", 4243 => "0000000000000000", 4244 => "0000000000000000", 4245 => "0000000000000000", 4246 => "0000000000000000", 4247 => "0000000000000000", 4248 => "0000000000000000", 4249 => "0000000000000000", 4250 => "0000000000000000", 4251 => "0000000000000000", 4252 => "0000000000000000", 4253 => "0000000000000000", 4254 => "0000000000000000", 4255 => "0000000000000000", 4256 => "0000000000000000", 4257 => "0000000000000000", 4258 => "0000000000000000", 4259 => "0000000000000000", 4260 => "0000000000000000", 4261 => "0000000000000000", 4262 => "0000000000000000", 4263 => "0000000000000000", 4264 => "0000000000000000", 4265 => "0000000000000000", 4266 => "0000000000000000", 4267 => "0000000000000000", 4268 => "0000000000000000", 4269 => "0000000000000000", 4270 => "0000000000000000", 4271 => "0000000000000000", 4272 => "0000000000000000", 4273 => "0000000000000000", 4274 => "0000000000000000", 4275 => "0000000000000000", 4276 => "0000000000000000", 4277 => "0000000000000000", 4278 => "0000000000000000", 4279 => "0000000000000000", 4280 => "0000000000000000", 4281 => "0000000000000000", 4282 => "0000000000000000", 4283 => "0000000000000000", 4284 => "0000000000000000", 4285 => "0000000000000000", 4286 => "0000000000000000", 4287 => "0000000000000000", 4288 => "0000000000000000", 4289 => "0000000000000000", 4290 => "0000000000000000", 4291 => "0000000000000000", 4292 => "0000000000000000", 4293 => "0000000000000000", 4294 => "0000000000000000", 4295 => "0000000000000000", 4296 => "0000000000000000", 4297 => "0000000000000000", 4298 => "0000000000000000", 4299 => "0000000000000000", 4300 => "0000000000000000", 4301 => "0000000000000000", 4302 => "0000000000000000", 4303 => "0000000000000000", 4304 => "0000000000000000", 4305 => "0000000000000000", 4306 => "0000000000000000", 4307 => "0000000000000000", 4308 => "0000000000000000", 4309 => "0000000000000000", 4310 => "0000000000000000", 4311 => "0000000000000000", 4312 => "0000000000000000", 4313 => "0000000000000000", 4314 => "0000000000000000", 4315 => "0000000000000000", 4316 => "0000000000000000", 4317 => "0000000000000000", 4318 => "0000000000000000", 4319 => "0000000000000000", 4320 => "0000000000000000", 4321 => "0000000000000000", 4322 => "0000000000000000", 4323 => "0000000000000000", 4324 => "0000000000000000", 4325 => "0000000000000000", 4326 => "0000000000000000", 4327 => "0000000000000000", 4328 => "0000000000000000", 4329 => "0000000000000000", 4330 => "0000000000000000", 4331 => "0000000000000000", 4332 => "0000000000000000", 4333 => "0000000000000000", 4334 => "0000000000000000", 4335 => "0000000000000000", 4336 => "0000000000000000", 4337 => "0000000000000000", 4338 => "0000000000000000", 4339 => "0000000000000000", 4340 => "0000000000000000", 4341 => "0000000000000000", 4342 => "0000000000000000", 4343 => "0000000000000000", 4344 => "0000000000000000", 4345 => "0000000000000000", 4346 => "0000000000000000", 4347 => "0000000000000000", 4348 => "0000000000000000", 4349 => "0000000000000000", 4350 => "0000000000000000", 4351 => "0000000000000000", 4352 => "0000000000000000", 4353 => "0000000000000000", 4354 => "0000000000000000", 4355 => "0000000000000000", 4356 => "0000000000000000", 4357 => "0000000000000000", 4358 => "0000000000000000", 4359 => "0000000000000000", 4360 => "0000000000000000", 4361 => "0000000000000000", 4362 => "0000000000000000", 4363 => "0000000000000000", 4364 => "0000000000000000", 4365 => "0000000000000000", 4366 => "0000000000000000", 4367 => "0000000000000000", 4368 => "0000000000000000", 4369 => "0000000000000000", 4370 => "0000000000000000", 4371 => "0000000000000000", 4372 => "0000000000000000", 4373 => "0000000000000000", 4374 => "0000000000000000", 4375 => "0000000000000000", 4376 => "0000000000000000", 4377 => "0000000000000000", 4378 => "0000000000000000", 4379 => "0000000000000000", 4380 => "0000000000000000", 4381 => "0000000000000000", 4382 => "0000000000000000", 4383 => "0000000000000000", 4384 => "0000000000000000", 4385 => "0000000000000000", 4386 => "0000000000000000", 4387 => "0000000000000000", 4388 => "0000000000000000", 4389 => "0000000000000000", 4390 => "0000000000000000", 4391 => "0000000000000000", 4392 => "0000000000000000", 4393 => "0000000000000000", 4394 => "0000000000000000", 4395 => "0000000000000000", 4396 => "0000000000000000", 4397 => "0000000000000000", 4398 => "0000000000000000", 4399 => "0000000000000000", 4400 => "0000000000000000", 4401 => "0000000000000000", 4402 => "0000000000000000", 4403 => "0000000000000000", 4404 => "0000000000000000", 4405 => "0000000000000000", 4406 => "0000000000000000", 4407 => "0000000000000000", 4408 => "0000000000000000", 4409 => "0000000000000000", 4410 => "0000000000000000", 4411 => "0000000000000000", 4412 => "0000000000000000", 4413 => "0000000000000000", 4414 => "0000000000000000", 4415 => "0000000000000000", 4416 => "0000000000000000", 4417 => "0000000000000000", 4418 => "0000000000000000", 4419 => "0000000000000000", 4420 => "0000000000000000", 4421 => "0000000000000000", 4422 => "0000000000000000", 4423 => "0000000000000000", 4424 => "0000000000000000", 4425 => "0000000000000000", 4426 => "0000000000000000", 4427 => "0000000000000000", 4428 => "0000000000000000", 4429 => "0000000000000000", 4430 => "0000000000000000", 4431 => "0000000000000000", 4432 => "0000000000000000", 4433 => "0000000000000000", 4434 => "0000000000000000", 4435 => "0000000000000000", 4436 => "0000000000000000", 4437 => "0000000000000000", 4438 => "0000000000000000", 4439 => "0000000000000000", 4440 => "0000000000000000", 4441 => "0000000000000000", 4442 => "0000000000000000", 4443 => "0000000000000000", 4444 => "0000000000000000", 4445 => "0000000000000000", 4446 => "0000000000000000", 4447 => "0000000000000000", 4448 => "0000000000000000", 4449 => "0000000000000000", 4450 => "0000000000000000", 4451 => "0000000000000000", 4452 => "0000000000000000", 4453 => "0000000000000000", 4454 => "0000000000000000", 4455 => "0000000000000000", 4456 => "0000000000000000", 4457 => "0000000000000000", 4458 => "0000000000000000", 4459 => "0000000000000000", 4460 => "0000000000000000", 4461 => "0000000000000000", 4462 => "0000000000000000", 4463 => "0000000000000000", 4464 => "0000000000000000", 4465 => "0000000000000000", 4466 => "0000000000000000", 4467 => "0000000000000000", 4468 => "0000000000000000", 4469 => "0000000000000000", 4470 => "0000000000000000", 4471 => "0000000000000000", 4472 => "0000000000000000", 4473 => "0000000000000000", 4474 => "0000000000000000", 4475 => "0000000000000000", 4476 => "0000000000000000", 4477 => "0000000000000000", 4478 => "0000000000000000", 4479 => "0000000000000000", 4480 => "0000000000000000", 4481 => "0000000000000000", 4482 => "0000000000000000", 4483 => "0000000000000000", 4484 => "0000000000000000", 4485 => "0000000000000000", 4486 => "0000000000000000", 4487 => "0000000000000000", 4488 => "0000000000000000", 4489 => "0000000000000000", 4490 => "0000000000000000", 4491 => "0000000000000000", 4492 => "0000000000000000", 4493 => "0000000000000000", 4494 => "0000000000000000", 4495 => "0000000000000000", 4496 => "0000000000000000", 4497 => "0000000000000000", 4498 => "0000000000000000", 4499 => "0000000000000000", 4500 => "0000000000000000", 4501 => "0000000000000000", 4502 => "0000000000000000", 4503 => "0000000000000000", 4504 => "0000000000000000", 4505 => "0000000000000000", 4506 => "0000000000000000", 4507 => "0000000000000000", 4508 => "0000000000000000", 4509 => "0000000000000000", 4510 => "0000000000000000", 4511 => "0000000000000000", 4512 => "0000000000000000", 4513 => "0000000000000000", 4514 => "0000000000000000", 4515 => "0000000000000000", 4516 => "0000000000000000", 4517 => "0000000000000000", 4518 => "0000000000000000", 4519 => "0000000000000000", 4520 => "0000000000000000", 4521 => "0000000000000000", 4522 => "0000000000000000", 4523 => "0000000000000000", 4524 => "0000000000000000", 4525 => "0000000000000000", 4526 => "0000000000000000", 4527 => "0000000000000000", 4528 => "0000000000000000", 4529 => "0000000000000000", 4530 => "0000000000000000", 4531 => "0000000000000000", 4532 => "0000000000000000", 4533 => "0000000000000000", 4534 => "0000000000000000", 4535 => "0000000000000000", 4536 => "0000000000000000", 4537 => "0000000000000000", 4538 => "0000000000000000", 4539 => "0000000000000000", 4540 => "0000000000000000", 4541 => "0000000000000000", 4542 => "0000000000000000", 4543 => "0000000000000000", 4544 => "0000000000000000", 4545 => "0000000000000000", 4546 => "0000000000000000", 4547 => "0000000000000000", 4548 => "0000000000000000", 4549 => "0000000000000000", 4550 => "0000000000000000", 4551 => "0000000000000000", 4552 => "0000000000000000", 4553 => "0000000000000000", 4554 => "0000000000000000", 4555 => "0000000000000000", 4556 => "0000000000000000", 4557 => "0000000000000000", 4558 => "0000000000000000", 4559 => "0000000000000000", 4560 => "0000000000000000", 4561 => "0000000000000000", 4562 => "0000000000000000", 4563 => "0000000000000000", 4564 => "0000000000000000", 4565 => "0000000000000000", 4566 => "0000000000000000", 4567 => "0000000000000000", 4568 => "0000000000000000", 4569 => "0000000000000000", 4570 => "0000000000000000", 4571 => "0000000000000000", 4572 => "0000000000000000", 4573 => "0000000000000000", 4574 => "0000000000000000", 4575 => "0000000000000000", 4576 => "0000000000000000", 4577 => "0000000000000000", 4578 => "0000000000000000", 4579 => "0000000000000000", 4580 => "0000000000000000", 4581 => "0000000000000000", 4582 => "0000000000000000", 4583 => "0000000000000000", 4584 => "0000000000000000", 4585 => "0000000000000000", 4586 => "0000000000000000", 4587 => "0000000000000000", 4588 => "0000000000000000", 4589 => "0000000000000000", 4590 => "0000000000000000", 4591 => "0000000000000000", 4592 => "0000000000000000", 4593 => "0000000000000000", 4594 => "0000000000000000", 4595 => "0000000000000000", 4596 => "0000000000000000", 4597 => "0000000000000000", 4598 => "0000000000000000", 4599 => "0000000000000000", 4600 => "0000000000000000", 4601 => "0000000000000000", 4602 => "0000000000000000", 4603 => "0000000000000000", 4604 => "0000000000000000", 4605 => "0000000000000000", 4606 => "0000000000000000", 4607 => "0000000000000000", 4608 => "0000000000000000", 4609 => "0000000000000000", 4610 => "0000000000000000", 4611 => "0000000000000000", 4612 => "0000000000000000", 4613 => "0000000000000000", 4614 => "0000000000000000", 4615 => "0000000000000000", 4616 => "0000000000000000", 4617 => "0000000000000000", 4618 => "0000000000000000", 4619 => "0000000000000000", 4620 => "0000000000000000", 4621 => "0000000000000000", 4622 => "0000000000000000", 4623 => "0000000000000000", 4624 => "0000000000000000", 4625 => "0000000000000000", 4626 => "0000000000000000", 4627 => "0000000000000000", 4628 => "0000000000000000", 4629 => "0000000000000000", 4630 => "0000000000000000", 4631 => "0000000000000000", 4632 => "0000000000000000", 4633 => "0000000000000000", 4634 => "0000000000000000", 4635 => "0000000000000000", 4636 => "0000000000000000", 4637 => "0000000000000000", 4638 => "0000000000000000", 4639 => "0000000000000000", 4640 => "0000000000000000", 4641 => "0000000000000000", 4642 => "0000000000000000", 4643 => "0000000000000000", 4644 => "0000000000000000", 4645 => "0000000000000000", 4646 => "0000000000000000", 4647 => "0000000000000000", 4648 => "0000000000000000", 4649 => "0000000000000000", 4650 => "0000000000000000", 4651 => "0000000000000000", 4652 => "0000000000000000", 4653 => "0000000000000000", 4654 => "0000000000000000", 4655 => "0000000000000000", 4656 => "0000000000000000", 4657 => "0000000000000000", 4658 => "0000000000000000", 4659 => "0000000000000000", 4660 => "0000000000000000", 4661 => "0000000000000000", 4662 => "0000000000000000", 4663 => "0000000000000000", 4664 => "0000000000000000", 4665 => "0000000000000000", 4666 => "0000000000000000", 4667 => "0000000000000000", 4668 => "0000000000000000", 4669 => "0000000000000000", 4670 => "0000000000000000", 4671 => "0000000000000000", 4672 => "0000000000000000", 4673 => "0000000000000000", 4674 => "0000000000000000", 4675 => "0000000000000000", 4676 => "0000000000000000", 4677 => "0000000000000000", 4678 => "0000000000000000", 4679 => "0000000000000000", 4680 => "0000000000000000", 4681 => "0000000000000000", 4682 => "0000000000000000", 4683 => "0000000000000000", 4684 => "0000000000000000", 4685 => "0000000000000000", 4686 => "0000000000000000", 4687 => "0000000000000000", 4688 => "0000000000000000", 4689 => "0000000000000000", 4690 => "0000000000000000", 4691 => "0000000000000000", 4692 => "0000000000000000", 4693 => "0000000000000000", 4694 => "0000000000000000", 4695 => "0000000000000000", 4696 => "0000000000000000", 4697 => "0000000000000000", 4698 => "0000000000000000", 4699 => "0000000000000000", 4700 => "0000000000000000", 4701 => "0000000000000000", 4702 => "0000000000000000", 4703 => "0000000000000000", 4704 => "0000000000000000", 4705 => "0000000000000000", 4706 => "0000000000000000", 4707 => "0000000000000000", 4708 => "0000000000000000", 4709 => "0000000000000000", 4710 => "0000000000000000", 4711 => "0000000000000000", 4712 => "0000000000000000", 4713 => "0000000000000000", 4714 => "0000000000000000", 4715 => "0000000000000000", 4716 => "0000000000000000", 4717 => "0000000000000000", 4718 => "0000000000000000", 4719 => "0000000000000000", 4720 => "0000000000000000", 4721 => "0000000000000000", 4722 => "0000000000000000", 4723 => "0000000000000000", 4724 => "0000000000000000", 4725 => "0000000000000000", 4726 => "0000000000000000", 4727 => "0000000000000000", 4728 => "0000000000000000", 4729 => "0000000000000000", 4730 => "0000000000000000", 4731 => "0000000000000000", 4732 => "0000000000000000", 4733 => "0000000000000000", 4734 => "0000000000000000", 4735 => "0000000000000000", 4736 => "0000000000000000", 4737 => "0000000000000000", 4738 => "0000000000000000", 4739 => "0000000000000000", 4740 => "0000000000000000", 4741 => "0000000000000000", 4742 => "0000000000000000", 4743 => "0000000000000000", 4744 => "0000000000000000", 4745 => "0000000000000000", 4746 => "0000000000000000", 4747 => "0000000000000000", 4748 => "0000000000000000", 4749 => "0000000000000000", 4750 => "0000000000000000", 4751 => "0000000000000000", 4752 => "0000000000000000", 4753 => "0000000000000000", 4754 => "0000000000000000", 4755 => "0000000000000000", 4756 => "0000000000000000", 4757 => "0000000000000000", 4758 => "0000000000000000", 4759 => "0000000000000000", 4760 => "0000000000000000", 4761 => "0000000000000000", 4762 => "0000000000000000", 4763 => "0000000000000000", 4764 => "0000000000000000", 4765 => "0000000000000000", 4766 => "0000000000000000", 4767 => "0000000000000000", 4768 => "0000000000000000", 4769 => "0000000000000000", 4770 => "0000000000000000", 4771 => "0000000000000000", 4772 => "0000000000000000", 4773 => "0000000000000000", 4774 => "0000000000000000", 4775 => "0000000000000000", 4776 => "0000000000000000", 4777 => "0000000000000000", 4778 => "0000000000000000", 4779 => "0000000000000000", 4780 => "0000000000000000", 4781 => "0000000000000000", 4782 => "0000000000000000", 4783 => "0000000000000000", 4784 => "0000000000000000", 4785 => "0000000000000000", 4786 => "0000000000000000", 4787 => "0000000000000000", 4788 => "0000000000000000", 4789 => "0000000000000000", 4790 => "0000000000000000", 4791 => "0000000000000000", 4792 => "0000000000000000", 4793 => "0000000000000000", 4794 => "0000000000000000", 4795 => "0000000000000000", 4796 => "0000000000000000", 4797 => "0000000000000000", 4798 => "0000000000000000", 4799 => "0000000000000000", 4800 => "0000000000000000", 4801 => "0000000000000000", 4802 => "0000000000000000", 4803 => "0000000000000000", 4804 => "0000000000000000", 4805 => "0000000000000000", 4806 => "0000000000000000", 4807 => "0000000000000000", 4808 => "0000000000000000", 4809 => "0000000000000000", 4810 => "0000000000000000", 4811 => "0000000000000000", 4812 => "0000000000000000", 4813 => "0000000000000000", 4814 => "0000000000000000", 4815 => "0000000000000000", 4816 => "0000000000000000", 4817 => "0000000000000000", 4818 => "0000000000000000", 4819 => "0000000000000000", 4820 => "0000000000000000", 4821 => "0000000000000000", 4822 => "0000000000000000", 4823 => "0000000000000000", 4824 => "0000000000000000", 4825 => "0000000000000000", 4826 => "0000000000000000", 4827 => "0000000000000000", 4828 => "0000000000000000", 4829 => "0000000000000000", 4830 => "0000000000000000", 4831 => "0000000000000000", 4832 => "0000000000000000", 4833 => "0000000000000000", 4834 => "0000000000000000", 4835 => "0000000000000000", 4836 => "0000000000000000", 4837 => "0000000000000000", 4838 => "0000000000000000", 4839 => "0000000000000000", 4840 => "0000000000000000", 4841 => "0000000000000000", 4842 => "0000000000000000", 4843 => "0000000000000000", 4844 => "0000000000000000", 4845 => "0000000000000000", 4846 => "0000000000000000", 4847 => "0000000000000000", 4848 => "0000000000000000", 4849 => "0000000000000000", 4850 => "0000000000000000", 4851 => "0000000000000000", 4852 => "0000000000000000", 4853 => "0000000000000000", 4854 => "0000000000000000", 4855 => "0000000000000000", 4856 => "0000000000000000", 4857 => "0000000000000000", 4858 => "0000000000000000", 4859 => "0000000000000000", 4860 => "0000000000000000", 4861 => "0000000000000000", 4862 => "0000000000000000", 4863 => "0000000000000000", 4864 => "0000000000000000", 4865 => "0000000000000000", 4866 => "0000000000000000", 4867 => "0000000000000000", 4868 => "0000000000000000", 4869 => "0000000000000000", 4870 => "0000000000000000", 4871 => "0000000000000000", 4872 => "0000000000000000", 4873 => "0000000000000000", 4874 => "0000000000000000", 4875 => "0000000000000000", 4876 => "0000000000000000", 4877 => "0000000000000000", 4878 => "0000000000000000", 4879 => "0000000000000000", 4880 => "0000000000000000", 4881 => "0000000000000000", 4882 => "0000000000000000", 4883 => "0000000000000000", 4884 => "0000000000000000", 4885 => "0000000000000000", 4886 => "0000000000000000", 4887 => "0000000000000000", 4888 => "0000000000000000", 4889 => "0000000000000000", 4890 => "0000000000000000", 4891 => "0000000000000000", 4892 => "0000000000000000", 4893 => "0000000000000000", 4894 => "0000000000000000", 4895 => "0000000000000000", 4896 => "0000000000000000", 4897 => "0000000000000000", 4898 => "0000000000000000", 4899 => "0000000000000000", 4900 => "0000000000000000", 4901 => "0000000000000000", 4902 => "0000000000000000", 4903 => "0000000000000000", 4904 => "0000000000000000", 4905 => "0000000000000000", 4906 => "0000000000000000", 4907 => "0000000000000000", 4908 => "0000000000000000", 4909 => "0000000000000000", 4910 => "0000000000000000", 4911 => "0000000000000000", 4912 => "0000000000000000", 4913 => "0000000000000000", 4914 => "0000000000000000", 4915 => "0000000000000000", 4916 => "0000000000000000", 4917 => "0000000000000000", 4918 => "0000000000000000", 4919 => "0000000000000000", 4920 => "0000000000000000", 4921 => "0000000000000000", 4922 => "0000000000000000", 4923 => "0000000000000000", 4924 => "0000000000000000", 4925 => "0000000000000000", 4926 => "0000000000000000", 4927 => "0000000000000000", 4928 => "0000000000000000", 4929 => "0000000000000000", 4930 => "0000000000000000", 4931 => "0000000000000000", 4932 => "0000000000000000", 4933 => "0000000000000000", 4934 => "0000000000000000", 4935 => "0000000000000000", 4936 => "0000000000000000", 4937 => "0000000000000000", 4938 => "0000000000000000", 4939 => "0000000000000000", 4940 => "0000000000000000", 4941 => "0000000000000000", 4942 => "0000000000000000", 4943 => "0000000000000000", 4944 => "0000000000000000", 4945 => "0000000000000000", 4946 => "0000000000000000", 4947 => "0000000000000000", 4948 => "0000000000000000", 4949 => "0000000000000000", 4950 => "0000000000000000", 4951 => "0000000000000000", 4952 => "0000000000000000", 4953 => "0000000000000000", 4954 => "0000000000000000", 4955 => "0000000000000000", 4956 => "0000000000000000", 4957 => "0000000000000000", 4958 => "0000000000000000", 4959 => "0000000000000000", 4960 => "0000000000000000", 4961 => "0000000000000000", 4962 => "0000000000000000", 4963 => "0000000000000000", 4964 => "0000000000000000", 4965 => "0000000000000000", 4966 => "0000000000000000", 4967 => "0000000000000000", 4968 => "0000000000000000", 4969 => "0000000000000000", 4970 => "0000000000000000", 4971 => "0000000000000000", 4972 => "0000000000000000", 4973 => "0000000000000000", 4974 => "0000000000000000", 4975 => "0000000000000000", 4976 => "0000000000000000", 4977 => "0000000000000000", 4978 => "0000000000000000", 4979 => "0000000000000000", 4980 => "0000000000000000", 4981 => "0000000000000000", 4982 => "0000000000000000", 4983 => "0000000000000000", 4984 => "0000000000000000", 4985 => "0000000000000000", 4986 => "0000000000000000", 4987 => "0000000000000000", 4988 => "0000000000000000", 4989 => "0000000000000000", 4990 => "0000000000000000", 4991 => "0000000000000000", 4992 => "0000000000000000", 4993 => "0000000000000000", 4994 => "0000000000000000", 4995 => "0000000000000000", 4996 => "0000000000000000", 4997 => "0000000000000000", 4998 => "0000000000000000", 4999 => "0000000000000000", 5000 => "0000000000000000", 5001 => "0000000000000000", 5002 => "0000000000000000", 5003 => "0000000000000000", 5004 => "0000000000000000", 5005 => "0000000000000000", 5006 => "0000000000000000", 5007 => "0000000000000000", 5008 => "0000000000000000", 5009 => "0000000000000000", 5010 => "0000000000000000", 5011 => "0000000000000000", 5012 => "0000000000000000", 5013 => "0000000000000000", 5014 => "0000000000000000", 5015 => "0000000000000000", 5016 => "0000000000000000", 5017 => "0000000000000000", 5018 => "0000000000000000", 5019 => "0000000000000000", 5020 => "0000000000000000", 5021 => "0000000000000000", 5022 => "0000000000000000", 5023 => "0000000000000000", 5024 => "0000000000000000", 5025 => "0000000000000000", 5026 => "0000000000000000", 5027 => "0000000000000000", 5028 => "0000000000000000", 5029 => "0000000000000000", 5030 => "0000000000000000", 5031 => "0000000000000000", 5032 => "0000000000000000", 5033 => "0000000000000000", 5034 => "0000000000000000", 5035 => "0000000000000000", 5036 => "0000000000000000", 5037 => "0000000000000000", 5038 => "0000000000000000", 5039 => "0000000000000000", 5040 => "0000000000000000", 5041 => "0000000000000000", 5042 => "0000000000000000", 5043 => "0000000000000000", 5044 => "0000000000000000", 5045 => "0000000000000000", 5046 => "0000000000000000", 5047 => "0000000000000000", 5048 => "0000000000000000", 5049 => "0000000000000000", 5050 => "0000000000000000", 5051 => "0000000000000000", 5052 => "0000000000000000", 5053 => "0000000000000000", 5054 => "0000000000000000", 5055 => "0000000000000000", 5056 => "0000000000000000", 5057 => "0000000000000000", 5058 => "0000000000000000", 5059 => "0000000000000000", 5060 => "0000000000000000", 5061 => "0000000000000000", 5062 => "0000000000000000", 5063 => "0000000000000000", 5064 => "0000000000000000", 5065 => "0000000000000000", 5066 => "0000000000000000", 5067 => "0000000000000000", 5068 => "0000000000000000", 5069 => "0000000000000000", 5070 => "0000000000000000", 5071 => "0000000000000000", 5072 => "0000000000000000", 5073 => "0000000000000000", 5074 => "0000000000000000", 5075 => "0000000000000000", 5076 => "0000000000000000", 5077 => "0000000000000000", 5078 => "0000000000000000", 5079 => "0000000000000000", 5080 => "0000000000000000", 5081 => "0000000000000000", 5082 => "0000000000000000", 5083 => "0000000000000000", 5084 => "0000000000000000", 5085 => "0000000000000000", 5086 => "0000000000000000", 5087 => "0000000000000000", 5088 => "0000000000000000", 5089 => "0000000000000000", 5090 => "0000000000000000", 5091 => "0000000000000000", 5092 => "0000000000000000", 5093 => "0000000000000000", 5094 => "0000000000000000", 5095 => "0000000000000000", 5096 => "0000000000000000", 5097 => "0000000000000000", 5098 => "0000000000000000", 5099 => "0000000000000000", 5100 => "0000000000000000", 5101 => "0000000000000000", 5102 => "0000000000000000", 5103 => "0000000000000000", 5104 => "0000000000000000", 5105 => "0000000000000000", 5106 => "0000000000000000", 5107 => "0000000000000000", 5108 => "0000000000000000", 5109 => "0000000000000000", 5110 => "0000000000000000", 5111 => "0000000000000000", 5112 => "0000000000000000", 5113 => "0000000000000000", 5114 => "0000000000000000", 5115 => "0000000000000000", 5116 => "0000000000000000", 5117 => "0000000000000000", 5118 => "0000000000000000", 5119 => "0000000000000000", 5120 => "0000000000000000", 5121 => "0000000000000000", 5122 => "0000000000000000", 5123 => "0000000000000000", 5124 => "0000000000000000", 5125 => "0000000000000000", 5126 => "0000000000000000", 5127 => "0000000000000000", 5128 => "0000000000000000", 5129 => "0000000000000000", 5130 => "0000000000000000", 5131 => "0000000000000000", 5132 => "0000000000000000", 5133 => "0000000000000000", 5134 => "0000000000000000", 5135 => "0000000000000000", 5136 => "0000000000000000", 5137 => "0000000000000000", 5138 => "0000000000000000", 5139 => "0000000000000000", 5140 => "0000000000000000", 5141 => "0000000000000000", 5142 => "0000000000000000", 5143 => "0000000000000000", 5144 => "0000000000000000", 5145 => "0000000000000000", 5146 => "0000000000000000", 5147 => "0000000000000000", 5148 => "0000000000000000", 5149 => "0000000000000000", 5150 => "0000000000000000", 5151 => "0000000000000000", 5152 => "0000000000000000", 5153 => "0000000000000000", 5154 => "0000000000000000", 5155 => "0000000000000000", 5156 => "0000000000000000", 5157 => "0000000000000000", 5158 => "0000000000000000", 5159 => "0000000000000000", 5160 => "0000000000000000", 5161 => "0000000000000000", 5162 => "0000000000000000", 5163 => "0000000000000000", 5164 => "0000000000000000", 5165 => "0000000000000000", 5166 => "0000000000000000", 5167 => "0000000000000000", 5168 => "0000000000000000", 5169 => "0000000000000000", 5170 => "0000000000000000", 5171 => "0000000000000000", 5172 => "0000000000000000", 5173 => "0000000000000000", 5174 => "0000000000000000", 5175 => "0000000000000000", 5176 => "0000000000000000", 5177 => "0000000000000000", 5178 => "0000000000000000", 5179 => "0000000000000000", 5180 => "0000000000000000", 5181 => "0000000000000000", 5182 => "0000000000000000", 5183 => "0000000000000000", 5184 => "0000000000000000", 5185 => "0000000000000000", 5186 => "0000000000000000", 5187 => "0000000000000000", 5188 => "0000000000000000", 5189 => "0000000000000000", 5190 => "0000000000000000", 5191 => "0000000000000000", 5192 => "0000000000000000", 5193 => "0000000000000000", 5194 => "0000000000000000", 5195 => "0000000000000000", 5196 => "0000000000000000", 5197 => "0000000000000000", 5198 => "0000000000000000", 5199 => "0000000000000000", 5200 => "0000000000000000", 5201 => "0000000000000000", 5202 => "0000000000000000", 5203 => "0000000000000000", 5204 => "0000000000000000", 5205 => "0000000000000000", 5206 => "0000000000000000", 5207 => "0000000000000000", 5208 => "0000000000000000", 5209 => "0000000000000000", 5210 => "0000000000000000", 5211 => "0000000000000000", 5212 => "0000000000000000", 5213 => "0000000000000000", 5214 => "0000000000000000", 5215 => "0000000000000000", 5216 => "0000000000000000", 5217 => "0000000000000000", 5218 => "0000000000000000", 5219 => "0000000000000000", 5220 => "0000000000000000", 5221 => "0000000000000000", 5222 => "0000000000000000", 5223 => "0000000000000000", 5224 => "0000000000000000", 5225 => "0000000000000000", 5226 => "0000000000000000", 5227 => "0000000000000000", 5228 => "0000000000000000", 5229 => "0000000000000000", 5230 => "0000000000000000", 5231 => "0000000000000000", 5232 => "0000000000000000", 5233 => "0000000000000000", 5234 => "0000000000000000", 5235 => "0000000000000000", 5236 => "0000000000000000", 5237 => "0000000000000000", 5238 => "0000000000000000", 5239 => "0000000000000000", 5240 => "0000000000000000", 5241 => "0000000000000000", 5242 => "0000000000000000", 5243 => "0000000000000000", 5244 => "0000000000000000", 5245 => "0000000000000000", 5246 => "0000000000000000", 5247 => "0000000000000000", 5248 => "0000000000000000", 5249 => "0000000000000000", 5250 => "0000000000000000", 5251 => "0000000000000000", 5252 => "0000000000000000", 5253 => "0000000000000000", 5254 => "0000000000000000", 5255 => "0000000000000000", 5256 => "0000000000000000", 5257 => "0000000000000000", 5258 => "0000000000000000", 5259 => "0000000000000000", 5260 => "0000000000000000", 5261 => "0000000000000000", 5262 => "0000000000000000", 5263 => "0000000000000000", 5264 => "0000000000000000", 5265 => "0000000000000000", 5266 => "0000000000000000", 5267 => "0000000000000000", 5268 => "0000000000000000", 5269 => "0000000000000000", 5270 => "0000000000000000", 5271 => "0000000000000000", 5272 => "0000000000000000", 5273 => "0000000000000000", 5274 => "0000000000000000", 5275 => "0000000000000000", 5276 => "0000000000000000", 5277 => "0000000000000000", 5278 => "0000000000000000", 5279 => "0000000000000000", 5280 => "0000000000000000", 5281 => "0000000000000000", 5282 => "0000000000000000", 5283 => "0000000000000000", 5284 => "0000000000000000", 5285 => "0000000000000000", 5286 => "0000000000000000", 5287 => "0000000000000000", 5288 => "0000000000000000", 5289 => "0000000000000000", 5290 => "0000000000000000", 5291 => "0000000000000000", 5292 => "0000000000000000", 5293 => "0000000000000000", 5294 => "0000000000000000", 5295 => "0000000000000000", 5296 => "0000000000000000", 5297 => "0000000000000000", 5298 => "0000000000000000", 5299 => "0000000000000000", 5300 => "0000000000000000", 5301 => "0000000000000000", 5302 => "0000000000000000", 5303 => "0000000000000000", 5304 => "0000000000000000", 5305 => "0000000000000000", 5306 => "0000000000000000", 5307 => "0000000000000000", 5308 => "0000000000000000", 5309 => "0000000000000000", 5310 => "0000000000000000", 5311 => "0000000000000000", 5312 => "0000000000000000", 5313 => "0000000000000000", 5314 => "0000000000000000", 5315 => "0000000000000000", 5316 => "0000000000000000", 5317 => "0000000000000000", 5318 => "0000000000000000", 5319 => "0000000000000000", 5320 => "0000000000000000", 5321 => "0000000000000000", 5322 => "0000000000000000", 5323 => "0000000000000000", 5324 => "0000000000000000", 5325 => "0000000000000000", 5326 => "0000000000000000", 5327 => "0000000000000000", 5328 => "0000000000000000", 5329 => "0000000000000000", 5330 => "0000000000000000", 5331 => "0000000000000000", 5332 => "0000000000000000", 5333 => "0000000000000000", 5334 => "0000000000000000", 5335 => "0000000000000000", 5336 => "0000000000000000", 5337 => "0000000000000000", 5338 => "0000000000000000", 5339 => "0000000000000000", 5340 => "0000000000000000", 5341 => "0000000000000000", 5342 => "0000000000000000", 5343 => "0000000000000000", 5344 => "0000000000000000", 5345 => "0000000000000000", 5346 => "0000000000000000", 5347 => "0000000000000000", 5348 => "0000000000000000", 5349 => "0000000000000000", 5350 => "0000000000000000", 5351 => "0000000000000000", 5352 => "0000000000000000", 5353 => "0000000000000000", 5354 => "0000000000000000", 5355 => "0000000000000000", 5356 => "0000000000000000", 5357 => "0000000000000000", 5358 => "0000000000000000", 5359 => "0000000000000000", 5360 => "0000000000000000", 5361 => "0000000000000000", 5362 => "0000000000000000", 5363 => "0000000000000000", 5364 => "0000000000000000", 5365 => "0000000000000000", 5366 => "0000000000000000", 5367 => "0000000000000000", 5368 => "0000000000000000", 5369 => "0000000000000000", 5370 => "0000000000000000", 5371 => "0000000000000000", 5372 => "0000000000000000", 5373 => "0000000000000000", 5374 => "0000000000000000", 5375 => "0000000000000000", 5376 => "0000000000000000", 5377 => "0000000000000000", 5378 => "0000000000000000", 5379 => "0000000000000000", 5380 => "0000000000000000", 5381 => "0000000000000000", 5382 => "0000000000000000", 5383 => "0000000000000000", 5384 => "0000000000000000", 5385 => "0000000000000000", 5386 => "0000000000000000", 5387 => "0000000000000000", 5388 => "0000000000000000", 5389 => "0000000000000000", 5390 => "0000000000000000", 5391 => "0000000000000000", 5392 => "0000000000000000", 5393 => "0000000000000000", 5394 => "0000000000000000", 5395 => "0000000000000000", 5396 => "0000000000000000", 5397 => "0000000000000000", 5398 => "0000000000000000", 5399 => "0000000000000000", 5400 => "0000000000000000", 5401 => "0000000000000000", 5402 => "0000000000000000", 5403 => "0000000000000000", 5404 => "0000000000000000", 5405 => "0000000000000000", 5406 => "0000000000000000", 5407 => "0000000000000000", 5408 => "0000000000000000", 5409 => "0000000000000000", 5410 => "0000000000000000", 5411 => "0000000000000000", 5412 => "0000000000000000", 5413 => "0000000000000000", 5414 => "0000000000000000", 5415 => "0000000000000000", 5416 => "0000000000000000", 5417 => "0000000000000000", 5418 => "0000000000000000", 5419 => "0000000000000000", 5420 => "0000000000000000", 5421 => "0000000000000000", 5422 => "0000000000000000", 5423 => "0000000000000000", 5424 => "0000000000000000", 5425 => "0000000000000000", 5426 => "0000000000000000", 5427 => "0000000000000000", 5428 => "0000000000000000", 5429 => "0000000000000000", 5430 => "0000000000000000", 5431 => "0000000000000000", 5432 => "0000000000000000", 5433 => "0000000000000000", 5434 => "0000000000000000", 5435 => "0000000000000000", 5436 => "0000000000000000", 5437 => "0000000000000000", 5438 => "0000000000000000", 5439 => "0000000000000000", 5440 => "0000000000000000", 5441 => "0000000000000000", 5442 => "0000000000000000", 5443 => "0000000000000000", 5444 => "0000000000000000", 5445 => "0000000000000000", 5446 => "0000000000000000", 5447 => "0000000000000000", 5448 => "0000000000000000", 5449 => "0000000000000000", 5450 => "0000000000000000", 5451 => "0000000000000000", 5452 => "0000000000000000", 5453 => "0000000000000000", 5454 => "0000000000000000", 5455 => "0000000000000000", 5456 => "0000000000000000", 5457 => "0000000000000000", 5458 => "0000000000000000", 5459 => "0000000000000000", 5460 => "0000000000000000", 5461 => "0000000000000000", 5462 => "0000000000000000", 5463 => "0000000000000000", 5464 => "0000000000000000", 5465 => "0000000000000000", 5466 => "0000000000000000", 5467 => "0000000000000000", 5468 => "0000000000000000", 5469 => "0000000000000000", 5470 => "0000000000000000", 5471 => "0000000000000000", 5472 => "0000000000000000", 5473 => "0000000000000000", 5474 => "0000000000000000", 5475 => "0000000000000000", 5476 => "0000000000000000", 5477 => "0000000000000000", 5478 => "0000000000000000", 5479 => "0000000000000000", 5480 => "0000000000000000", 5481 => "0000000000000000", 5482 => "0000000000000000", 5483 => "0000000000000000", 5484 => "0000000000000000", 5485 => "0000000000000000", 5486 => "0000000000000000", 5487 => "0000000000000000", 5488 => "0000000000000000", 5489 => "0000000000000000", 5490 => "0000000000000000", 5491 => "0000000000000000", 5492 => "0000000000000000", 5493 => "0000000000000000", 5494 => "0000000000000000", 5495 => "0000000000000000", 5496 => "0000000000000000", 5497 => "0000000000000000", 5498 => "0000000000000000", 5499 => "0000000000000000", 5500 => "0000000000000000", 5501 => "0000000000000000", 5502 => "0000000000000000", 5503 => "0000000000000000", 5504 => "0000000000000000", 5505 => "0000000000000000", 5506 => "0000000000000000", 5507 => "0000000000000000", 5508 => "0000000000000000", 5509 => "0000000000000000", 5510 => "0000000000000000", 5511 => "0000000000000000", 5512 => "0000000000000000", 5513 => "0000000000000000", 5514 => "0000000000000000", 5515 => "0000000000000000", 5516 => "0000000000000000", 5517 => "0000000000000000", 5518 => "0000000000000000", 5519 => "0000000000000000", 5520 => "0000000000000000", 5521 => "0000000000000000", 5522 => "0000000000000000", 5523 => "0000000000000000", 5524 => "0000000000000000", 5525 => "0000000000000000", 5526 => "0000000000000000", 5527 => "0000000000000000", 5528 => "0000000000000000", 5529 => "0000000000000000", 5530 => "0000000000000000", 5531 => "0000000000000000", 5532 => "0000000000000000", 5533 => "0000000000000000", 5534 => "0000000000000000", 5535 => "0000000000000000", 5536 => "0000000000000000", 5537 => "0000000000000000", 5538 => "0000000000000000", 5539 => "0000000000000000", 5540 => "0000000000000000", 5541 => "0000000000000000", 5542 => "0000000000000000", 5543 => "0000000000000000", 5544 => "0000000000000000", 5545 => "0000000000000000", 5546 => "0000000000000000", 5547 => "0000000000000000", 5548 => "0000000000000000", 5549 => "0000000000000000", 5550 => "0000000000000000", 5551 => "0000000000000000", 5552 => "0000000000000000", 5553 => "0000000000000000", 5554 => "0000000000000000", 5555 => "0000000000000000", 5556 => "0000000000000000", 5557 => "0000000000000000", 5558 => "0000000000000000", 5559 => "0000000000000000", 5560 => "0000000000000000", 5561 => "0000000000000000", 5562 => "0000000000000000", 5563 => "0000000000000000", 5564 => "0000000000000000", 5565 => "0000000000000000", 5566 => "0000000000000000", 5567 => "0000000000000000", 5568 => "0000000000000000", 5569 => "0000000000000000", 5570 => "0000000000000000", 5571 => "0000000000000000", 5572 => "0000000000000000", 5573 => "0000000000000000", 5574 => "0000000000000000", 5575 => "0000000000000000", 5576 => "0000000000000000", 5577 => "0000000000000000", 5578 => "0000000000000000", 5579 => "0000000000000000", 5580 => "0000000000000000", 5581 => "0000000000000000", 5582 => "0000000000000000", 5583 => "0000000000000000", 5584 => "0000000000000000", 5585 => "0000000000000000", 5586 => "0000000000000000", 5587 => "0000000000000000", 5588 => "0000000000000000", 5589 => "0000000000000000", 5590 => "0000000000000000", 5591 => "0000000000000000", 5592 => "0000000000000000", 5593 => "0000000000000000", 5594 => "0000000000000000", 5595 => "0000000000000000", 5596 => "0000000000000000", 5597 => "0000000000000000", 5598 => "0000000000000000", 5599 => "0000000000000000", 5600 => "0000000000000000", 5601 => "0000000000000000", 5602 => "0000000000000000", 5603 => "0000000000000000", 5604 => "0000000000000000", 5605 => "0000000000000000", 5606 => "0000000000000000", 5607 => "0000000000000000", 5608 => "0000000000000000", 5609 => "0000000000000000", 5610 => "0000000000000000", 5611 => "0000000000000000", 5612 => "0000000000000000", 5613 => "0000000000000000", 5614 => "0000000000000000", 5615 => "0000000000000000", 5616 => "0000000000000000", 5617 => "0000000000000000", 5618 => "0000000000000000", 5619 => "0000000000000000", 5620 => "0000000000000000", 5621 => "0000000000000000", 5622 => "0000000000000000", 5623 => "0000000000000000", 5624 => "0000000000000000", 5625 => "0000000000000000", 5626 => "0000000000000000", 5627 => "0000000000000000", 5628 => "0000000000000000", 5629 => "0000000000000000", 5630 => "0000000000000000", 5631 => "0000000000000000", 5632 => "0000000000000000", 5633 => "0000000000000000", 5634 => "0000000000000000", 5635 => "0000000000000000", 5636 => "0000000000000000", 5637 => "0000000000000000", 5638 => "0000000000000000", 5639 => "0000000000000000", 5640 => "0000000000000000", 5641 => "0000000000000000", 5642 => "0000000000000000", 5643 => "0000000000000000", 5644 => "0000000000000000", 5645 => "0000000000000000", 5646 => "0000000000000000", 5647 => "0000000000000000", 5648 => "0000000000000000", 5649 => "0000000000000000", 5650 => "0000000000000000", 5651 => "0000000000000000", 5652 => "0000000000000000", 5653 => "0000000000000000", 5654 => "0000000000000000", 5655 => "0000000000000000", 5656 => "0000000000000000", 5657 => "0000000000000000", 5658 => "0000000000000000", 5659 => "0000000000000000", 5660 => "0000000000000000", 5661 => "0000000000000000", 5662 => "0000000000000000", 5663 => "0000000000000000", 5664 => "0000000000000000", 5665 => "0000000000000000", 5666 => "0000000000000000", 5667 => "0000000000000000", 5668 => "0000000000000000", 5669 => "0000000000000000", 5670 => "0000000000000000", 5671 => "0000000000000000", 5672 => "0000000000000000", 5673 => "0000000000000000", 5674 => "0000000000000000", 5675 => "0000000000000000", 5676 => "0000000000000000", 5677 => "0000000000000000", 5678 => "0000000000000000", 5679 => "0000000000000000", 5680 => "0000000000000000", 5681 => "0000000000000000", 5682 => "0000000000000000", 5683 => "0000000000000000", 5684 => "0000000000000000", 5685 => "0000000000000000", 5686 => "0000000000000000", 5687 => "0000000000000000", 5688 => "0000000000000000", 5689 => "0000000000000000", 5690 => "0000000000000000", 5691 => "0000000000000000", 5692 => "0000000000000000", 5693 => "0000000000000000", 5694 => "0000000000000000", 5695 => "0000000000000000", 5696 => "0000000000000000", 5697 => "0000000000000000", 5698 => "0000000000000000", 5699 => "0000000000000000", 5700 => "0000000000000000", 5701 => "0000000000000000", 5702 => "0000000000000000", 5703 => "0000000000000000", 5704 => "0000000000000000", 5705 => "0000000000000000", 5706 => "0000000000000000", 5707 => "0000000000000000", 5708 => "0000000000000000", 5709 => "0000000000000000", 5710 => "0000000000000000", 5711 => "0000000000000000", 5712 => "0000000000000000", 5713 => "0000000000000000", 5714 => "0000000000000000", 5715 => "0000000000000000", 5716 => "0000000000000000", 5717 => "0000000000000000", 5718 => "0000000000000000", 5719 => "0000000000000000", 5720 => "0000000000000000", 5721 => "0000000000000000", 5722 => "0000000000000000", 5723 => "0000000000000000", 5724 => "0000000000000000", 5725 => "0000000000000000", 5726 => "0000000000000000", 5727 => "0000000000000000", 5728 => "0000000000000000", 5729 => "0000000000000000", 5730 => "0000000000000000", 5731 => "0000000000000000", 5732 => "0000000000000000", 5733 => "0000000000000000", 5734 => "0000000000000000", 5735 => "0000000000000000", 5736 => "0000000000000000", 5737 => "0000000000000000", 5738 => "0000000000000000", 5739 => "0000000000000000", 5740 => "0000000000000000", 5741 => "0000000000000000", 5742 => "0000000000000000", 5743 => "0000000000000000", 5744 => "0000000000000000", 5745 => "0000000000000000", 5746 => "0000000000000000", 5747 => "0000000000000000", 5748 => "0000000000000000", 5749 => "0000000000000000", 5750 => "0000000000000000", 5751 => "0000000000000000", 5752 => "0000000000000000", 5753 => "0000000000000000", 5754 => "0000000000000000", 5755 => "0000000000000000", 5756 => "0000000000000000", 5757 => "0000000000000000", 5758 => "0000000000000000", 5759 => "0000000000000000", 5760 => "0000000000000000", 5761 => "0000000000000000", 5762 => "0000000000000000", 5763 => "0000000000000000", 5764 => "0000000000000000", 5765 => "0000000000000000", 5766 => "0000000000000000", 5767 => "0000000000000000", 5768 => "0000000000000000", 5769 => "0000000000000000", 5770 => "0000000000000000", 5771 => "0000000000000000", 5772 => "0000000000000000", 5773 => "0000000000000000", 5774 => "0000000000000000", 5775 => "0000000000000000", 5776 => "0000000000000000", 5777 => "0000000000000000", 5778 => "0000000000000000", 5779 => "0000000000000000", 5780 => "0000000000000000", 5781 => "0000000000000000", 5782 => "0000000000000000", 5783 => "0000000000000000", 5784 => "0000000000000000", 5785 => "0000000000000000", 5786 => "0000000000000000", 5787 => "0000000000000000", 5788 => "0000000000000000", 5789 => "0000000000000000", 5790 => "0000000000000000", 5791 => "0000000000000000", 5792 => "0000000000000000", 5793 => "0000000000000000", 5794 => "0000000000000000", 5795 => "0000000000000000", 5796 => "0000000000000000", 5797 => "0000000000000000", 5798 => "0000000000000000", 5799 => "0000000000000000", 5800 => "0000000000000000", 5801 => "0000000000000000", 5802 => "0000000000000000", 5803 => "0000000000000000", 5804 => "0000000000000000", 5805 => "0000000000000000", 5806 => "0000000000000000", 5807 => "0000000000000000", 5808 => "0000000000000000", 5809 => "0000000000000000", 5810 => "0000000000000000", 5811 => "0000000000000000", 5812 => "0000000000000000", 5813 => "0000000000000000", 5814 => "0000000000000000", 5815 => "0000000000000000", 5816 => "0000000000000000", 5817 => "0000000000000000", 5818 => "0000000000000000", 5819 => "0000000000000000", 5820 => "0000000000000000", 5821 => "0000000000000000", 5822 => "0000000000000000", 5823 => "0000000000000000", 5824 => "0000000000000000", 5825 => "0000000000000000", 5826 => "0000000000000000", 5827 => "0000000000000000", 5828 => "0000000000000000", 5829 => "0000000000000000", 5830 => "0000000000000000", 5831 => "0000000000000000", 5832 => "0000000000000000", 5833 => "0000000000000000", 5834 => "0000000000000000", 5835 => "0000000000000000", 5836 => "0000000000000000", 5837 => "0000000000000000", 5838 => "0000000000000000", 5839 => "0000000000000000", 5840 => "0000000000000000", 5841 => "0000000000000000", 5842 => "0000000000000000", 5843 => "0000000000000000", 5844 => "0000000000000000", 5845 => "0000000000000000", 5846 => "0000000000000000", 5847 => "0000000000000000", 5848 => "0000000000000000", 5849 => "0000000000000000", 5850 => "0000000000000000", 5851 => "0000000000000000", 5852 => "0000000000000000", 5853 => "0000000000000000", 5854 => "0000000000000000", 5855 => "0000000000000000", 5856 => "0000000000000000", 5857 => "0000000000000000", 5858 => "0000000000000000", 5859 => "0000000000000000", 5860 => "0000000000000000", 5861 => "0000000000000000", 5862 => "0000000000000000", 5863 => "0000000000000000", 5864 => "0000000000000000", 5865 => "0000000000000000", 5866 => "0000000000000000", 5867 => "0000000000000000", 5868 => "0000000000000000", 5869 => "0000000000000000", 5870 => "0000000000000000", 5871 => "0000000000000000", 5872 => "0000000000000000", 5873 => "0000000000000000", 5874 => "0000000000000000", 5875 => "0000000000000000", 5876 => "0000000000000000", 5877 => "0000000000000000", 5878 => "0000000000000000", 5879 => "0000000000000000", 5880 => "0000000000000000", 5881 => "0000000000000000", 5882 => "0000000000000000", 5883 => "0000000000000000", 5884 => "0000000000000000", 5885 => "0000000000000000", 5886 => "0000000000000000", 5887 => "0000000000000000", 5888 => "0000000000000000", 5889 => "0000000000000000", 5890 => "0000000000000000", 5891 => "0000000000000000", 5892 => "0000000000000000", 5893 => "0000000000000000", 5894 => "0000000000000000", 5895 => "0000000000000000", 5896 => "0000000000000000", 5897 => "0000000000000000", 5898 => "0000000000000000", 5899 => "0000000000000000", 5900 => "0000000000000000", 5901 => "0000000000000000", 5902 => "0000000000000000", 5903 => "0000000000000000", 5904 => "0000000000000000", 5905 => "0000000000000000", 5906 => "0000000000000000", 5907 => "0000000000000000", 5908 => "0000000000000000", 5909 => "0000000000000000", 5910 => "0000000000000000", 5911 => "0000000000000000", 5912 => "0000000000000000", 5913 => "0000000000000000", 5914 => "0000000000000000", 5915 => "0000000000000000", 5916 => "0000000000000000", 5917 => "0000000000000000", 5918 => "0000000000000000", 5919 => "0000000000000000", 5920 => "0000000000000000", 5921 => "0000000000000000", 5922 => "0000000000000000", 5923 => "0000000000000000", 5924 => "0000000000000000", 5925 => "0000000000000000", 5926 => "0000000000000000", 5927 => "0000000000000000", 5928 => "0000000000000000", 5929 => "0000000000000000", 5930 => "0000000000000000", 5931 => "0000000000000000", 5932 => "0000000000000000", 5933 => "0000000000000000", 5934 => "0000000000000000", 5935 => "0000000000000000", 5936 => "0000000000000000", 5937 => "0000000000000000", 5938 => "0000000000000000", 5939 => "0000000000000000", 5940 => "0000000000000000", 5941 => "0000000000000000", 5942 => "0000000000000000", 5943 => "0000000000000000", 5944 => "0000000000000000", 5945 => "0000000000000000", 5946 => "0000000000000000", 5947 => "0000000000000000", 5948 => "0000000000000000", 5949 => "0000000000000000", 5950 => "0000000000000000", 5951 => "0000000000000000", 5952 => "0000000000000000", 5953 => "0000000000000000", 5954 => "0000000000000000", 5955 => "0000000000000000", 5956 => "0000000000000000", 5957 => "0000000000000000", 5958 => "0000000000000000", 5959 => "0000000000000000", 5960 => "0000000000000000", 5961 => "0000000000000000", 5962 => "0000000000000000", 5963 => "0000000000000000", 5964 => "0000000000000000", 5965 => "0000000000000000", 5966 => "0000000000000000", 5967 => "0000000000000000", 5968 => "0000000000000000", 5969 => "0000000000000000", 5970 => "0000000000000000", 5971 => "0000000000000000", 5972 => "0000000000000000", 5973 => "0000000000000000", 5974 => "0000000000000000", 5975 => "0000000000000000", 5976 => "0000000000000000", 5977 => "0000000000000000", 5978 => "0000000000000000", 5979 => "0000000000000000", 5980 => "0000000000000000", 5981 => "0000000000000000", 5982 => "0000000000000000", 5983 => "0000000000000000", 5984 => "0000000000000000", 5985 => "0000000000000000", 5986 => "0000000000000000", 5987 => "0000000000000000", 5988 => "0000000000000000", 5989 => "0000000000000000", 5990 => "0000000000000000", 5991 => "0000000000000000", 5992 => "0000000000000000", 5993 => "0000000000000000", 5994 => "0000000000000000", 5995 => "0000000000000000", 5996 => "0000000000000000", 5997 => "0000000000000000", 5998 => "0000000000000000", 5999 => "0000000000000000", 6000 => "0000000000000000", 6001 => "0000000000000000", 6002 => "0000000000000000", 6003 => "0000000000000000", 6004 => "0000000000000000", 6005 => "0000000000000000", 6006 => "0000000000000000", 6007 => "0000000000000000", 6008 => "0000000000000000", 6009 => "0000000000000000", 6010 => "0000000000000000", 6011 => "0000000000000000", 6012 => "0000000000000000", 6013 => "0000000000000000", 6014 => "0000000000000000", 6015 => "0000000000000000", 6016 => "0000000000000000", 6017 => "0000000000000000", 6018 => "0000000000000000", 6019 => "0000000000000000", 6020 => "0000000000000000", 6021 => "0000000000000000", 6022 => "0000000000000000", 6023 => "0000000000000000", 6024 => "0000000000000000", 6025 => "0000000000000000", 6026 => "0000000000000000", 6027 => "0000000000000000", 6028 => "0000000000000000", 6029 => "0000000000000000", 6030 => "0000000000000000", 6031 => "0000000000000000", 6032 => "0000000000000000", 6033 => "0000000000000000", 6034 => "0000000000000000", 6035 => "0000000000000000", 6036 => "0000000000000000", 6037 => "0000000000000000", 6038 => "0000000000000000", 6039 => "0000000000000000", 6040 => "0000000000000000", 6041 => "0000000000000000", 6042 => "0000000000000000", 6043 => "0000000000000000", 6044 => "0000000000000000", 6045 => "0000000000000000", 6046 => "0000000000000000", 6047 => "0000000000000000", 6048 => "0000000000000000", 6049 => "0000000000000000", 6050 => "0000000000000000", 6051 => "0000000000000000", 6052 => "0000000000000000", 6053 => "0000000000000000", 6054 => "0000000000000000", 6055 => "0000000000000000", 6056 => "0000000000000000", 6057 => "0000000000000000", 6058 => "0000000000000000", 6059 => "0000000000000000", 6060 => "0000000000000000", 6061 => "0000000000000000", 6062 => "0000000000000000", 6063 => "0000000000000000", 6064 => "0000000000000000", 6065 => "0000000000000000", 6066 => "0000000000000000", 6067 => "0000000000000000", 6068 => "0000000000000000", 6069 => "0000000000000000", 6070 => "0000000000000000", 6071 => "0000000000000000", 6072 => "0000000000000000", 6073 => "0000000000000000", 6074 => "0000000000000000", 6075 => "0000000000000000", 6076 => "0000000000000000", 6077 => "0000000000000000", 6078 => "0000000000000000", 6079 => "0000000000000000", 6080 => "0000000000000000", 6081 => "0000000000000000", 6082 => "0000000000000000", 6083 => "0000000000000000", 6084 => "0000000000000000", 6085 => "0000000000000000", 6086 => "0000000000000000", 6087 => "0000000000000000", 6088 => "0000000000000000", 6089 => "0000000000000000", 6090 => "0000000000000000", 6091 => "0000000000000000", 6092 => "0000000000000000", 6093 => "0000000000000000", 6094 => "0000000000000000", 6095 => "0000000000000000", 6096 => "0000000000000000", 6097 => "0000000000000000", 6098 => "0000000000000000", 6099 => "0000000000000000", 6100 => "0000000000000000", 6101 => "0000000000000000", 6102 => "0000000000000000", 6103 => "0000000000000000", 6104 => "0000000000000000", 6105 => "0000000000000000", 6106 => "0000000000000000", 6107 => "0000000000000000", 6108 => "0000000000000000", 6109 => "0000000000000000", 6110 => "0000000000000000", 6111 => "0000000000000000", 6112 => "0000000000000000", 6113 => "0000000000000000", 6114 => "0000000000000000", 6115 => "0000000000000000", 6116 => "0000000000000000", 6117 => "0000000000000000", 6118 => "0000000000000000", 6119 => "0000000000000000", 6120 => "0000000000000000", 6121 => "0000000000000000", 6122 => "0000000000000000", 6123 => "0000000000000000", 6124 => "0000000000000000", 6125 => "0000000000000000", 6126 => "0000000000000000", 6127 => "0000000000000000", 6128 => "0000000000000000", 6129 => "0000000000000000", 6130 => "0000000000000000", 6131 => "0000000000000000", 6132 => "0000000000000000", 6133 => "0000000000000000", 6134 => "0000000000000000", 6135 => "0000000000000000", 6136 => "0000000000000000", 6137 => "0000000000000000", 6138 => "0000000000000000", 6139 => "0000000000000000", 6140 => "0000000000000000", 6141 => "0000000000000000", 6142 => "0000000000000000", 6143 => "0000000000000000", 6144 => "0000000000000000", 6145 => "0000000000000000", 6146 => "0000000000000000", 6147 => "0000000000000000", 6148 => "0000000000000000", 6149 => "0000000000000000", 6150 => "0000000000000000", 6151 => "0000000000000000", 6152 => "0000000000000000", 6153 => "0000000000000000", 6154 => "0000000000000000", 6155 => "0000000000000000", 6156 => "0000000000000000", 6157 => "0000000000000000", 6158 => "0000000000000000", 6159 => "0000000000000000", 6160 => "0000000000000000", 6161 => "0000000000000000", 6162 => "0000000000000000", 6163 => "0000000000000000", 6164 => "0000000000000000", 6165 => "0000000000000000", 6166 => "0000000000000000", 6167 => "0000000000000000", 6168 => "0000000000000000", 6169 => "0000000000000000", 6170 => "0000000000000000", 6171 => "0000000000000000", 6172 => "0000000000000000", 6173 => "0000000000000000", 6174 => "0000000000000000", 6175 => "0000000000000000", 6176 => "0000000000000000", 6177 => "0000000000000000", 6178 => "0000000000000000", 6179 => "0000000000000000", 6180 => "0000000000000000", 6181 => "0000000000000000", 6182 => "0000000000000000", 6183 => "0000000000000000", 6184 => "0000000000000000", 6185 => "0000000000000000", 6186 => "0000000000000000", 6187 => "0000000000000000", 6188 => "0000000000000000", 6189 => "0000000000000000", 6190 => "0000000000000000", 6191 => "0000000000000000", 6192 => "0000000000000000", 6193 => "0000000000000000", 6194 => "0000000000000000", 6195 => "0000000000000000", 6196 => "0000000000000000", 6197 => "0000000000000000", 6198 => "0000000000000000", 6199 => "0000000000000000", 6200 => "0000000000000000", 6201 => "0000000000000000", 6202 => "0000000000000000", 6203 => "0000000000000000", 6204 => "0000000000000000", 6205 => "0000000000000000", 6206 => "0000000000000000", 6207 => "0000000000000000", 6208 => "0000000000000000", 6209 => "0000000000000000", 6210 => "0000000000000000", 6211 => "0000000000000000", 6212 => "0000000000000000", 6213 => "0000000000000000", 6214 => "0000000000000000", 6215 => "0000000000000000", 6216 => "0000000000000000", 6217 => "0000000000000000", 6218 => "0000000000000000", 6219 => "0000000000000000", 6220 => "0000000000000000", 6221 => "0000000000000000", 6222 => "0000000000000000", 6223 => "0000000000000000", 6224 => "0000000000000000", 6225 => "0000000000000000", 6226 => "0000000000000000", 6227 => "0000000000000000", 6228 => "0000000000000000", 6229 => "0000000000000000", 6230 => "0000000000000000", 6231 => "0000000000000000", 6232 => "0000000000000000", 6233 => "0000000000000000", 6234 => "0000000000000000", 6235 => "0000000000000000", 6236 => "0000000000000000", 6237 => "0000000000000000", 6238 => "0000000000000000", 6239 => "0000000000000000", 6240 => "0000000000000000", 6241 => "0000000000000000", 6242 => "0000000000000000", 6243 => "0000000000000000", 6244 => "0000000000000000", 6245 => "0000000000000000", 6246 => "0000000000000000", 6247 => "0000000000000000", 6248 => "0000000000000000", 6249 => "0000000000000000", 6250 => "0000000000000000", 6251 => "0000000000000000", 6252 => "0000000000000000", 6253 => "0000000000000000", 6254 => "0000000000000000", 6255 => "0000000000000000", 6256 => "0000000000000000", 6257 => "0000000000000000", 6258 => "0000000000000000", 6259 => "0000000000000000", 6260 => "0000000000000000", 6261 => "0000000000000000", 6262 => "0000000000000000", 6263 => "0000000000000000", 6264 => "0000000000000000", 6265 => "0000000000000000", 6266 => "0000000000000000", 6267 => "0000000000000000", 6268 => "0000000000000000", 6269 => "0000000000000000", 6270 => "0000000000000000", 6271 => "0000000000000000", 6272 => "0000000000000000", 6273 => "0000000000000000", 6274 => "0000000000000000", 6275 => "0000000000000000", 6276 => "0000000000000000", 6277 => "0000000000000000", 6278 => "0000000000000000", 6279 => "0000000000000000", 6280 => "0000000000000000", 6281 => "0000000000000000", 6282 => "0000000000000000", 6283 => "0000000000000000", 6284 => "0000000000000000", 6285 => "0000000000000000", 6286 => "0000000000000000", 6287 => "0000000000000000", 6288 => "0000000000000000", 6289 => "0000000000000000", 6290 => "0000000000000000", 6291 => "0000000000000000", 6292 => "0000000000000000", 6293 => "0000000000000000", 6294 => "0000000000000000", 6295 => "0000000000000000", 6296 => "0000000000000000", 6297 => "0000000000000000", 6298 => "0000000000000000", 6299 => "0000000000000000", 6300 => "0000000000000000", 6301 => "0000000000000000", 6302 => "0000000000000000", 6303 => "0000000000000000", 6304 => "0000000000000000", 6305 => "0000000000000000", 6306 => "0000000000000000", 6307 => "0000000000000000", 6308 => "0000000000000000", 6309 => "0000000000000000", 6310 => "0000000000000000", 6311 => "0000000000000000", 6312 => "0000000000000000", 6313 => "0000000000000000", 6314 => "0000000000000000", 6315 => "0000000000000000", 6316 => "0000000000000000", 6317 => "0000000000000000", 6318 => "0000000000000000", 6319 => "0000000000000000", 6320 => "0000000000000000", 6321 => "0000000000000000", 6322 => "0000000000000000", 6323 => "0000000000000000", 6324 => "0000000000000000", 6325 => "0000000000000000", 6326 => "0000000000000000", 6327 => "0000000000000000", 6328 => "0000000000000000", 6329 => "0000000000000000", 6330 => "0000000000000000", 6331 => "0000000000000000", 6332 => "0000000000000000", 6333 => "0000000000000000", 6334 => "0000000000000000", 6335 => "0000000000000000", 6336 => "0000000000000000", 6337 => "0000000000000000", 6338 => "0000000000000000", 6339 => "0000000000000000", 6340 => "0000000000000000", 6341 => "0000000000000000", 6342 => "0000000000000000", 6343 => "0000000000000000", 6344 => "0000000000000000", 6345 => "0000000000000000", 6346 => "0000000000000000", 6347 => "0000000000000000", 6348 => "0000000000000000", 6349 => "0000000000000000", 6350 => "0000000000000000", 6351 => "0000000000000000", 6352 => "0000000000000000", 6353 => "0000000000000000", 6354 => "0000000000000000", 6355 => "0000000000000000", 6356 => "0000000000000000", 6357 => "0000000000000000", 6358 => "0000000000000000", 6359 => "0000000000000000", 6360 => "0000000000000000", 6361 => "0000000000000000", 6362 => "0000000000000000", 6363 => "0000000000000000", 6364 => "0000000000000000", 6365 => "0000000000000000", 6366 => "0000000000000000", 6367 => "0000000000000000", 6368 => "0000000000000000", 6369 => "0000000000000000", 6370 => "0000000000000000", 6371 => "0000000000000000", 6372 => "0000000000000000", 6373 => "0000000000000000", 6374 => "0000000000000000", 6375 => "0000000000000000", 6376 => "0000000000000000", 6377 => "0000000000000000", 6378 => "0000000000000000", 6379 => "0000000000000000", 6380 => "0000000000000000", 6381 => "0000000000000000", 6382 => "0000000000000000", 6383 => "0000000000000000", 6384 => "0000000000000000", 6385 => "0000000000000000", 6386 => "0000000000000000", 6387 => "0000000000000000", 6388 => "0000000000000000", 6389 => "0000000000000000", 6390 => "0000000000000000", 6391 => "0000000000000000", 6392 => "0000000000000000", 6393 => "0000000000000000", 6394 => "0000000000000000", 6395 => "0000000000000000", 6396 => "0000000000000000", 6397 => "0000000000000000", 6398 => "0000000000000000", 6399 => "0000000000000000", 6400 => "0000000000000000", 6401 => "0000000000000000", 6402 => "0000000000000000", 6403 => "0000000000000000", 6404 => "0000000000000000", 6405 => "0000000000000000", 6406 => "0000000000000000", 6407 => "0000000000000000", 6408 => "0000000000000000", 6409 => "0000000000000000", 6410 => "0000000000000000", 6411 => "0000000000000000", 6412 => "0000000000000000", 6413 => "0000000000000000", 6414 => "0000000000000000", 6415 => "0000000000000000", 6416 => "0000000000000000", 6417 => "0000000000000000", 6418 => "0000000000000000", 6419 => "0000000000000000", 6420 => "0000000000000000", 6421 => "0000000000000000", 6422 => "0000000000000000", 6423 => "0000000000000000", 6424 => "0000000000000000", 6425 => "0000000000000000", 6426 => "0000000000000000", 6427 => "0000000000000000", 6428 => "0000000000000000", 6429 => "0000000000000000", 6430 => "0000000000000000", 6431 => "0000000000000000", 6432 => "0000000000000000", 6433 => "0000000000000000", 6434 => "0000000000000000", 6435 => "0000000000000000", 6436 => "0000000000000000", 6437 => "0000000000000000", 6438 => "0000000000000000", 6439 => "0000000000000000", 6440 => "0000000000000000", 6441 => "0000000000000000", 6442 => "0000000000000000", 6443 => "0000000000000000", 6444 => "0000000000000000", 6445 => "0000000000000000", 6446 => "0000000000000000", 6447 => "0000000000000000", 6448 => "0000000000000000", 6449 => "0000000000000000", 6450 => "0000000000000000", 6451 => "0000000000000000", 6452 => "0000000000000000", 6453 => "0000000000000000", 6454 => "0000000000000000", 6455 => "0000000000000000", 6456 => "0000000000000000", 6457 => "0000000000000000", 6458 => "0000000000000000", 6459 => "0000000000000000", 6460 => "0000000000000000", 6461 => "0000000000000000", 6462 => "0000000000000000", 6463 => "0000000000000000", 6464 => "0000000000000000", 6465 => "0000000000000000", 6466 => "0000000000000000", 6467 => "0000000000000000", 6468 => "0000000000000000", 6469 => "0000000000000000", 6470 => "0000000000000000", 6471 => "0000000000000000", 6472 => "0000000000000000", 6473 => "0000000000000000", 6474 => "0000000000000000", 6475 => "0000000000000000", 6476 => "0000000000000000", 6477 => "0000000000000000", 6478 => "0000000000000000", 6479 => "0000000000000000", 6480 => "0000000000000000", 6481 => "0000000000000000", 6482 => "0000000000000000", 6483 => "0000000000000000", 6484 => "0000000000000000", 6485 => "0000000000000000", 6486 => "0000000000000000", 6487 => "0000000000000000", 6488 => "0000000000000000", 6489 => "0000000000000000", 6490 => "0000000000000000", 6491 => "0000000000000000", 6492 => "0000000000000000", 6493 => "0000000000000000", 6494 => "0000000000000000", 6495 => "0000000000000000", 6496 => "0000000000000000", 6497 => "0000000000000000", 6498 => "0000000000000000", 6499 => "0000000000000000", 6500 => "0000000000000000", 6501 => "0000000000000000", 6502 => "0000000000000000", 6503 => "0000000000000000", 6504 => "0000000000000000", 6505 => "0000000000000000", 6506 => "0000000000000000", 6507 => "0000000000000000", 6508 => "0000000000000000", 6509 => "0000000000000000", 6510 => "0000000000000000", 6511 => "0000000000000000", 6512 => "0000000000000000", 6513 => "0000000000000000", 6514 => "0000000000000000", 6515 => "0000000000000000", 6516 => "0000000000000000", 6517 => "0000000000000000", 6518 => "0000000000000000", 6519 => "0000000000000000", 6520 => "0000000000000000", 6521 => "0000000000000000", 6522 => "0000000000000000", 6523 => "0000000000000000", 6524 => "0000000000000000", 6525 => "0000000000000000", 6526 => "0000000000000000", 6527 => "0000000000000000", 6528 => "0000000000000000", 6529 => "0000000000000000", 6530 => "0000000000000000", 6531 => "0000000000000000", 6532 => "0000000000000000", 6533 => "0000000000000000", 6534 => "0000000000000000", 6535 => "0000000000000000", 6536 => "0000000000000000", 6537 => "0000000000000000", 6538 => "0000000000000000", 6539 => "0000000000000000", 6540 => "0000000000000000", 6541 => "0000000000000000", 6542 => "0000000000000000", 6543 => "0000000000000000", 6544 => "0000000000000000", 6545 => "0000000000000000", 6546 => "0000000000000000", 6547 => "0000000000000000", 6548 => "0000000000000000", 6549 => "0000000000000000", 6550 => "0000000000000000", 6551 => "0000000000000000", 6552 => "0000000000000000", 6553 => "0000000000000000", 6554 => "0000000000000000", 6555 => "0000000000000000", 6556 => "0000000000000000", 6557 => "0000000000000000", 6558 => "0000000000000000", 6559 => "0000000000000000", 6560 => "0000000000000000", 6561 => "0000000000000000", 6562 => "0000000000000000", 6563 => "0000000000000000", 6564 => "0000000000000000", 6565 => "0000000000000000", 6566 => "0000000000000000", 6567 => "0000000000000000", 6568 => "0000000000000000", 6569 => "0000000000000000", 6570 => "0000000000000000", 6571 => "0000000000000000", 6572 => "0000000000000000", 6573 => "0000000000000000", 6574 => "0000000000000000", 6575 => "0000000000000000", 6576 => "0000000000000000", 6577 => "0000000000000000", 6578 => "0000000000000000", 6579 => "0000000000000000", 6580 => "0000000000000000", 6581 => "0000000000000000", 6582 => "0000000000000000", 6583 => "0000000000000000", 6584 => "0000000000000000", 6585 => "0000000000000000", 6586 => "0000000000000000", 6587 => "0000000000000000", 6588 => "0000000000000000", 6589 => "0000000000000000", 6590 => "0000000000000000", 6591 => "0000000000000000", 6592 => "0000000000000000", 6593 => "0000000000000000", 6594 => "0000000000000000", 6595 => "0000000000000000", 6596 => "0000000000000000", 6597 => "0000000000000000", 6598 => "0000000000000000", 6599 => "0000000000000000", 6600 => "0000000000000000", 6601 => "0000000000000000", 6602 => "0000000000000000", 6603 => "0000000000000000", 6604 => "0000000000000000", 6605 => "0000000000000000", 6606 => "0000000000000000", 6607 => "0000000000000000", 6608 => "0000000000000000", 6609 => "0000000000000000", 6610 => "0000000000000000", 6611 => "0000000000000000", 6612 => "0000000000000000", 6613 => "0000000000000000", 6614 => "0000000000000000", 6615 => "0000000000000000", 6616 => "0000000000000000", 6617 => "0000000000000000", 6618 => "0000000000000000", 6619 => "0000000000000000", 6620 => "0000000000000000", 6621 => "0000000000000000", 6622 => "0000000000000000", 6623 => "0000000000000000", 6624 => "0000000000000000", 6625 => "0000000000000000", 6626 => "0000000000000000", 6627 => "0000000000000000", 6628 => "0000000000000000", 6629 => "0000000000000000", 6630 => "0000000000000000", 6631 => "0000000000000000", 6632 => "0000000000000000", 6633 => "0000000000000000", 6634 => "0000000000000000", 6635 => "0000000000000000", 6636 => "0000000000000000", 6637 => "0000000000000000", 6638 => "0000000000000000", 6639 => "0000000000000000", 6640 => "0000000000000000", 6641 => "0000000000000000", 6642 => "0000000000000000", 6643 => "0000000000000000", 6644 => "0000000000000000", 6645 => "0000000000000000", 6646 => "0000000000000000", 6647 => "0000000000000000", 6648 => "0000000000000000", 6649 => "0000000000000000", 6650 => "0000000000000000", 6651 => "0000000000000000", 6652 => "0000000000000000", 6653 => "0000000000000000", 6654 => "0000000000000000", 6655 => "0000000000000000", 6656 => "0000000000000000", 6657 => "0000000000000000", 6658 => "0000000000000000", 6659 => "0000000000000000", 6660 => "0000000000000000", 6661 => "0000000000000000", 6662 => "0000000000000000", 6663 => "0000000000000000", 6664 => "0000000000000000", 6665 => "0000000000000000", 6666 => "0000000000000000", 6667 => "0000000000000000", 6668 => "0000000000000000", 6669 => "0000000000000000", 6670 => "0000000000000000", 6671 => "0000000000000000", 6672 => "0000000000000000", 6673 => "0000000000000000", 6674 => "0000000000000000", 6675 => "0000000000000000", 6676 => "0000000000000000", 6677 => "0000000000000000", 6678 => "0000000000000000", 6679 => "0000000000000000", 6680 => "0000000000000000", 6681 => "0000000000000000", 6682 => "0000000000000000", 6683 => "0000000000000000", 6684 => "0000000000000000", 6685 => "0000000000000000", 6686 => "0000000000000000", 6687 => "0000000000000000", 6688 => "0000000000000000", 6689 => "0000000000000000", 6690 => "0000000000000000", 6691 => "0000000000000000", 6692 => "0000000000000000", 6693 => "0000000000000000", 6694 => "0000000000000000", 6695 => "0000000000000000", 6696 => "0000000000000000", 6697 => "0000000000000000", 6698 => "0000000000000000", 6699 => "0000000000000000", 6700 => "0000000000000000", 6701 => "0000000000000000", 6702 => "0000000000000000", 6703 => "0000000000000000", 6704 => "0000000000000000", 6705 => "0000000000000000", 6706 => "0000000000000000", 6707 => "0000000000000000", 6708 => "0000000000000000", 6709 => "0000000000000000", 6710 => "0000000000000000", 6711 => "0000000000000000", 6712 => "0000000000000000", 6713 => "0000000000000000", 6714 => "0000000000000000", 6715 => "0000000000000000", 6716 => "0000000000000000", 6717 => "0000000000000000", 6718 => "0000000000000000", 6719 => "0000000000000000", 6720 => "0000000000000000", 6721 => "0000000000000000", 6722 => "0000000000000000", 6723 => "0000000000000000", 6724 => "0000000000000000", 6725 => "0000000000000000", 6726 => "0000000000000000", 6727 => "0000000000000000", 6728 => "0000000000000000", 6729 => "0000000000000000", 6730 => "0000000000000000", 6731 => "0000000000000000", 6732 => "0000000000000000", 6733 => "0000000000000000", 6734 => "0000000000000000", 6735 => "0000000000000000", 6736 => "0000000000000000", 6737 => "0000000000000000", 6738 => "0000000000000000", 6739 => "0000000000000000", 6740 => "0000000000000000", 6741 => "0000000000000000", 6742 => "0000000000000000", 6743 => "0000000000000000", 6744 => "0000000000000000", 6745 => "0000000000000000", 6746 => "0000000000000000", 6747 => "0000000000000000", 6748 => "0000000000000000", 6749 => "0000000000000000", 6750 => "0000000000000000", 6751 => "0000000000000000", 6752 => "0000000000000000", 6753 => "0000000000000000", 6754 => "0000000000000000", 6755 => "0000000000000000", 6756 => "0000000000000000", 6757 => "0000000000000000", 6758 => "0000000000000000", 6759 => "0000000000000000", 6760 => "0000000000000000", 6761 => "0000000000000000", 6762 => "0000000000000000", 6763 => "0000000000000000", 6764 => "0000000000000000", 6765 => "0000000000000000", 6766 => "0000000000000000", 6767 => "0000000000000000", 6768 => "0000000000000000", 6769 => "0000000000000000", 6770 => "0000000000000000", 6771 => "0000000000000000", 6772 => "0000000000000000", 6773 => "0000000000000000", 6774 => "0000000000000000", 6775 => "0000000000000000", 6776 => "0000000000000000", 6777 => "0000000000000000", 6778 => "0000000000000000", 6779 => "0000000000000000", 6780 => "0000000000000000", 6781 => "0000000000000000", 6782 => "0000000000000000", 6783 => "0000000000000000", 6784 => "0000000000000000", 6785 => "0000000000000000", 6786 => "0000000000000000", 6787 => "0000000000000000", 6788 => "0000000000000000", 6789 => "0000000000000000", 6790 => "0000000000000000", 6791 => "0000000000000000", 6792 => "0000000000000000", 6793 => "0000000000000000", 6794 => "0000000000000000", 6795 => "0000000000000000", 6796 => "0000000000000000", 6797 => "0000000000000000", 6798 => "0000000000000000", 6799 => "0000000000000000", 6800 => "0000000000000000", 6801 => "0000000000000000", 6802 => "0000000000000000", 6803 => "0000000000000000", 6804 => "0000000000000000", 6805 => "0000000000000000", 6806 => "0000000000000000", 6807 => "0000000000000000", 6808 => "0000000000000000", 6809 => "0000000000000000", 6810 => "0000000000000000", 6811 => "0000000000000000", 6812 => "0000000000000000", 6813 => "0000000000000000", 6814 => "0000000000000000", 6815 => "0000000000000000", 6816 => "0000000000000000", 6817 => "0000000000000000", 6818 => "0000000000000000", 6819 => "0000000000000000", 6820 => "0000000000000000", 6821 => "0000000000000000", 6822 => "0000000000000000", 6823 => "0000000000000000", 6824 => "0000000000000000", 6825 => "0000000000000000", 6826 => "0000000000000000", 6827 => "0000000000000000", 6828 => "0000000000000000", 6829 => "0000000000000000", 6830 => "0000000000000000", 6831 => "0000000000000000", 6832 => "0000000000000000", 6833 => "0000000000000000", 6834 => "0000000000000000", 6835 => "0000000000000000", 6836 => "0000000000000000", 6837 => "0000000000000000", 6838 => "0000000000000000", 6839 => "0000000000000000", 6840 => "0000000000000000", 6841 => "0000000000000000", 6842 => "0000000000000000", 6843 => "0000000000000000", 6844 => "0000000000000000", 6845 => "0000000000000000", 6846 => "0000000000000000", 6847 => "0000000000000000", 6848 => "0000000000000000", 6849 => "0000000000000000", 6850 => "0000000000000000", 6851 => "0000000000000000", 6852 => "0000000000000000", 6853 => "0000000000000000", 6854 => "0000000000000000", 6855 => "0000000000000000", 6856 => "0000000000000000", 6857 => "0000000000000000", 6858 => "0000000000000000", 6859 => "0000000000000000", 6860 => "0000000000000000", 6861 => "0000000000000000", 6862 => "0000000000000000", 6863 => "0000000000000000", 6864 => "0000000000000000", 6865 => "0000000000000000", 6866 => "0000000000000000", 6867 => "0000000000000000", 6868 => "0000000000000000", 6869 => "0000000000000000", 6870 => "0000000000000000", 6871 => "0000000000000000", 6872 => "0000000000000000", 6873 => "0000000000000000", 6874 => "0000000000000000", 6875 => "0000000000000000", 6876 => "0000000000000000", 6877 => "0000000000000000", 6878 => "0000000000000000", 6879 => "0000000000000000", 6880 => "0000000000000000", 6881 => "0000000000000000", 6882 => "0000000000000000", 6883 => "0000000000000000", 6884 => "0000000000000000", 6885 => "0000000000000000", 6886 => "0000000000000000", 6887 => "0000000000000000", 6888 => "0000000000000000", 6889 => "0000000000000000", 6890 => "0000000000000000", 6891 => "0000000000000000", 6892 => "0000000000000000", 6893 => "0000000000000000", 6894 => "0000000000000000", 6895 => "0000000000000000", 6896 => "0000000000000000", 6897 => "0000000000000000", 6898 => "0000000000000000", 6899 => "0000000000000000", 6900 => "0000000000000000", 6901 => "0000000000000000", 6902 => "0000000000000000", 6903 => "0000000000000000", 6904 => "0000000000000000", 6905 => "0000000000000000", 6906 => "0000000000000000", 6907 => "0000000000000000", 6908 => "0000000000000000", 6909 => "0000000000000000", 6910 => "0000000000000000", 6911 => "0000000000000000", 6912 => "0000000000000000", 6913 => "0000000000000000", 6914 => "0000000000000000", 6915 => "0000000000000000", 6916 => "0000000000000000", 6917 => "0000000000000000", 6918 => "0000000000000000", 6919 => "0000000000000000", 6920 => "0000000000000000", 6921 => "0000000000000000", 6922 => "0000000000000000", 6923 => "0000000000000000", 6924 => "0000000000000000", 6925 => "0000000000000000", 6926 => "0000000000000000", 6927 => "0000000000000000", 6928 => "0000000000000000", 6929 => "0000000000000000", 6930 => "0000000000000000", 6931 => "0000000000000000", 6932 => "0000000000000000", 6933 => "0000000000000000", 6934 => "0000000000000000", 6935 => "0000000000000000", 6936 => "0000000000000000", 6937 => "0000000000000000", 6938 => "0000000000000000", 6939 => "0000000000000000", 6940 => "0000000000000000", 6941 => "0000000000000000", 6942 => "0000000000000000", 6943 => "0000000000000000", 6944 => "0000000000000000", 6945 => "0000000000000000", 6946 => "0000000000000000", 6947 => "0000000000000000", 6948 => "0000000000000000", 6949 => "0000000000000000", 6950 => "0000000000000000", 6951 => "0000000000000000", 6952 => "0000000000000000", 6953 => "0000000000000000", 6954 => "0000000000000000", 6955 => "0000000000000000", 6956 => "0000000000000000", 6957 => "0000000000000000", 6958 => "0000000000000000", 6959 => "0000000000000000", 6960 => "0000000000000000", 6961 => "0000000000000000", 6962 => "0000000000000000", 6963 => "0000000000000000", 6964 => "0000000000000000", 6965 => "0000000000000000", 6966 => "0000000000000000", 6967 => "0000000000000000", 6968 => "0000000000000000", 6969 => "0000000000000000", 6970 => "0000000000000000", 6971 => "0000000000000000", 6972 => "0000000000000000", 6973 => "0000000000000000", 6974 => "0000000000000000", 6975 => "0000000000000000", 6976 => "0000000000000000", 6977 => "0000000000000000", 6978 => "0000000000000000", 6979 => "0000000000000000", 6980 => "0000000000000000", 6981 => "0000000000000000", 6982 => "0000000000000000", 6983 => "0000000000000000", 6984 => "0000000000000000", 6985 => "0000000000000000", 6986 => "0000000000000000", 6987 => "0000000000000000", 6988 => "0000000000000000", 6989 => "0000000000000000", 6990 => "0000000000000000", 6991 => "0000000000000000", 6992 => "0000000000000000", 6993 => "0000000000000000", 6994 => "0000000000000000", 6995 => "0000000000000000", 6996 => "0000000000000000", 6997 => "0000000000000000", 6998 => "0000000000000000", 6999 => "0000000000000000", 7000 => "0000000000000000", 7001 => "0000000000000000", 7002 => "0000000000000000", 7003 => "0000000000000000", 7004 => "0000000000000000", 7005 => "0000000000000000", 7006 => "0000000000000000", 7007 => "0000000000000000", 7008 => "0000000000000000", 7009 => "0000000000000000", 7010 => "0000000000000000", 7011 => "0000000000000000", 7012 => "0000000000000000", 7013 => "0000000000000000", 7014 => "0000000000000000", 7015 => "0000000000000000", 7016 => "0000000000000000", 7017 => "0000000000000000", 7018 => "0000000000000000", 7019 => "0000000000000000", 7020 => "0000000000000000", 7021 => "0000000000000000", 7022 => "0000000000000000", 7023 => "0000000000000000", 7024 => "0000000000000000", 7025 => "0000000000000000", 7026 => "0000000000000000", 7027 => "0000000000000000", 7028 => "0000000000000000", 7029 => "0000000000000000", 7030 => "0000000000000000", 7031 => "0000000000000000", 7032 => "0000000000000000", 7033 => "0000000000000000", 7034 => "0000000000000000", 7035 => "0000000000000000", 7036 => "0000000000000000", 7037 => "0000000000000000", 7038 => "0000000000000000", 7039 => "0000000000000000", 7040 => "0000000000000000", 7041 => "0000000000000000", 7042 => "0000000000000000", 7043 => "0000000000000000", 7044 => "0000000000000000", 7045 => "0000000000000000", 7046 => "0000000000000000", 7047 => "0000000000000000", 7048 => "0000000000000000", 7049 => "0000000000000000", 7050 => "0000000000000000", 7051 => "0000000000000000", 7052 => "0000000000000000", 7053 => "0000000000000000", 7054 => "0000000000000000", 7055 => "0000000000000000", 7056 => "0000000000000000", 7057 => "0000000000000000", 7058 => "0000000000000000", 7059 => "0000000000000000", 7060 => "0000000000000000", 7061 => "0000000000000000", 7062 => "0000000000000000", 7063 => "0000000000000000", 7064 => "0000000000000000", 7065 => "0000000000000000", 7066 => "0000000000000000", 7067 => "0000000000000000", 7068 => "0000000000000000", 7069 => "0000000000000000", 7070 => "0000000000000000", 7071 => "0000000000000000", 7072 => "0000000000000000", 7073 => "0000000000000000", 7074 => "0000000000000000", 7075 => "0000000000000000", 7076 => "0000000000000000", 7077 => "0000000000000000", 7078 => "0000000000000000", 7079 => "0000000000000000", 7080 => "0000000000000000", 7081 => "0000000000000000", 7082 => "0000000000000000", 7083 => "0000000000000000", 7084 => "0000000000000000", 7085 => "0000000000000000", 7086 => "0000000000000000", 7087 => "0000000000000000", 7088 => "0000000000000000", 7089 => "0000000000000000", 7090 => "0000000000000000", 7091 => "0000000000000000", 7092 => "0000000000000000", 7093 => "0000000000000000", 7094 => "0000000000000000", 7095 => "0000000000000000", 7096 => "0000000000000000", 7097 => "0000000000000000", 7098 => "0000000000000000", 7099 => "0000000000000000", 7100 => "0000000000000000", 7101 => "0000000000000000", 7102 => "0000000000000000", 7103 => "0000000000000000", 7104 => "0000000000000000", 7105 => "0000000000000000", 7106 => "0000000000000000", 7107 => "0000000000000000", 7108 => "0000000000000000", 7109 => "0000000000000000", 7110 => "0000000000000000", 7111 => "0000000000000000", 7112 => "0000000000000000", 7113 => "0000000000000000", 7114 => "0000000000000000", 7115 => "0000000000000000", 7116 => "0000000000000000", 7117 => "0000000000000000", 7118 => "0000000000000000", 7119 => "0000000000000000", 7120 => "0000000000000000", 7121 => "0000000000000000", 7122 => "0000000000000000", 7123 => "0000000000000000", 7124 => "0000000000000000", 7125 => "0000000000000000", 7126 => "0000000000000000", 7127 => "0000000000000000", 7128 => "0000000000000000", 7129 => "0000000000000000", 7130 => "0000000000000000", 7131 => "0000000000000000", 7132 => "0000000000000000", 7133 => "0000000000000000", 7134 => "0000000000000000", 7135 => "0000000000000000", 7136 => "0000000000000000", 7137 => "0000000000000000", 7138 => "0000000000000000", 7139 => "0000000000000000", 7140 => "0000000000000000", 7141 => "0000000000000000", 7142 => "0000000000000000", 7143 => "0000000000000000", 7144 => "0000000000000000", 7145 => "0000000000000000", 7146 => "0000000000000000", 7147 => "0000000000000000", 7148 => "0000000000000000", 7149 => "0000000000000000", 7150 => "0000000000000000", 7151 => "0000000000000000", 7152 => "0000000000000000", 7153 => "0000000000000000", 7154 => "0000000000000000", 7155 => "0000000000000000", 7156 => "0000000000000000", 7157 => "0000000000000000", 7158 => "0000000000000000", 7159 => "0000000000000000", 7160 => "0000000000000000", 7161 => "0000000000000000", 7162 => "0000000000000000", 7163 => "0000000000000000", 7164 => "0000000000000000", 7165 => "0000000000000000", 7166 => "0000000000000000", 7167 => "0000000000000000", 7168 => "0000000000000000", 7169 => "0000000000000000", 7170 => "0000000000000000", 7171 => "0000000000000000", 7172 => "0000000000000000", 7173 => "0000000000000000", 7174 => "0000000000000000", 7175 => "0000000000000000", 7176 => "0000000000000000", 7177 => "0000000000000000", 7178 => "0000000000000000", 7179 => "0000000000000000", 7180 => "0000000000000000", 7181 => "0000000000000000", 7182 => "0000000000000000", 7183 => "0000000000000000", 7184 => "0000000000000000", 7185 => "0000000000000000", 7186 => "0000000000000000", 7187 => "0000000000000000", 7188 => "0000000000000000", 7189 => "0000000000000000", 7190 => "0000000000000000", 7191 => "0000000000000000", 7192 => "0000000000000000", 7193 => "0000000000000000", 7194 => "0000000000000000", 7195 => "0000000000000000", 7196 => "0000000000000000", 7197 => "0000000000000000", 7198 => "0000000000000000", 7199 => "0000000000000000", 7200 => "0000000000000000", 7201 => "0000000000000000", 7202 => "0000000000000000", 7203 => "0000000000000000", 7204 => "0000000000000000", 7205 => "0000000000000000", 7206 => "0000000000000000", 7207 => "0000000000000000", 7208 => "0000000000000000", 7209 => "0000000000000000", 7210 => "0000000000000000", 7211 => "0000000000000000", 7212 => "0000000000000000", 7213 => "0000000000000000", 7214 => "0000000000000000", 7215 => "0000000000000000", 7216 => "0000000000000000", 7217 => "0000000000000000", 7218 => "0000000000000000", 7219 => "0000000000000000", 7220 => "0000000000000000", 7221 => "0000000000000000", 7222 => "0000000000000000", 7223 => "0000000000000000", 7224 => "0000000000000000", 7225 => "0000000000000000", 7226 => "0000000000000000", 7227 => "0000000000000000", 7228 => "0000000000000000", 7229 => "0000000000000000", 7230 => "0000000000000000", 7231 => "0000000000000000", 7232 => "0000000000000000", 7233 => "0000000000000000", 7234 => "0000000000000000", 7235 => "0000000000000000", 7236 => "0000000000000000", 7237 => "0000000000000000", 7238 => "0000000000000000", 7239 => "0000000000000000", 7240 => "0000000000000000", 7241 => "0000000000000000", 7242 => "0000000000000000", 7243 => "0000000000000000", 7244 => "0000000000000000", 7245 => "0000000000000000", 7246 => "0000000000000000", 7247 => "0000000000000000", 7248 => "0000000000000000", 7249 => "0000000000000000", 7250 => "0000000000000000", 7251 => "0000000000000000", 7252 => "0000000000000000", 7253 => "0000000000000000", 7254 => "0000000000000000", 7255 => "0000000000000000", 7256 => "0000000000000000", 7257 => "0000000000000000", 7258 => "0000000000000000", 7259 => "0000000000000000", 7260 => "0000000000000000", 7261 => "0000000000000000", 7262 => "0000000000000000", 7263 => "0000000000000000", 7264 => "0000000000000000", 7265 => "0000000000000000", 7266 => "0000000000000000", 7267 => "0000000000000000", 7268 => "0000000000000000", 7269 => "0000000000000000", 7270 => "0000000000000000", 7271 => "0000000000000000", 7272 => "0000000000000000", 7273 => "0000000000000000", 7274 => "0000000000000000", 7275 => "0000000000000000", 7276 => "0000000000000000", 7277 => "0000000000000000", 7278 => "0000000000000000", 7279 => "0000000000000000", 7280 => "0000000000000000", 7281 => "0000000000000000", 7282 => "0000000000000000", 7283 => "0000000000000000", 7284 => "0000000000000000", 7285 => "0000000000000000", 7286 => "0000000000000000", 7287 => "0000000000000000", 7288 => "0000000000000000", 7289 => "0000000000000000", 7290 => "0000000000000000", 7291 => "0000000000000000", 7292 => "0000000000000000", 7293 => "0000000000000000", 7294 => "0000000000000000", 7295 => "0000000000000000", 7296 => "0000000000000000", 7297 => "0000000000000000", 7298 => "0000000000000000", 7299 => "0000000000000000", 7300 => "0000000000000000", 7301 => "0000000000000000", 7302 => "0000000000000000", 7303 => "0000000000000000", 7304 => "0000000000000000", 7305 => "0000000000000000", 7306 => "0000000000000000", 7307 => "0000000000000000", 7308 => "0000000000000000", 7309 => "0000000000000000", 7310 => "0000000000000000", 7311 => "0000000000000000", 7312 => "0000000000000000", 7313 => "0000000000000000", 7314 => "0000000000000000", 7315 => "0000000000000000", 7316 => "0000000000000000", 7317 => "0000000000000000", 7318 => "0000000000000000", 7319 => "0000000000000000", 7320 => "0000000000000000", 7321 => "0000000000000000", 7322 => "0000000000000000", 7323 => "0000000000000000", 7324 => "0000000000000000", 7325 => "0000000000000000", 7326 => "0000000000000000", 7327 => "0000000000000000", 7328 => "0000000000000000", 7329 => "0000000000000000", 7330 => "0000000000000000", 7331 => "0000000000000000", 7332 => "0000000000000000", 7333 => "0000000000000000", 7334 => "0000000000000000", 7335 => "0000000000000000", 7336 => "0000000000000000", 7337 => "0000000000000000", 7338 => "0000000000000000", 7339 => "0000000000000000", 7340 => "0000000000000000", 7341 => "0000000000000000", 7342 => "0000000000000000", 7343 => "0000000000000000", 7344 => "0000000000000000", 7345 => "0000000000000000", 7346 => "0000000000000000", 7347 => "0000000000000000", 7348 => "0000000000000000", 7349 => "0000000000000000", 7350 => "0000000000000000", 7351 => "0000000000000000", 7352 => "0000000000000000", 7353 => "0000000000000000", 7354 => "0000000000000000", 7355 => "0000000000000000", 7356 => "0000000000000000", 7357 => "0000000000000000", 7358 => "0000000000000000", 7359 => "0000000000000000", 7360 => "0000000000000000", 7361 => "0000000000000000", 7362 => "0000000000000000", 7363 => "0000000000000000", 7364 => "0000000000000000", 7365 => "0000000000000000", 7366 => "0000000000000000", 7367 => "0000000000000000", 7368 => "0000000000000000", 7369 => "0000000000000000", 7370 => "0000000000000000", 7371 => "0000000000000000", 7372 => "0000000000000000", 7373 => "0000000000000000", 7374 => "0000000000000000", 7375 => "0000000000000000", 7376 => "0000000000000000", 7377 => "0000000000000000", 7378 => "0000000000000000", 7379 => "0000000000000000", 7380 => "0000000000000000", 7381 => "0000000000000000", 7382 => "0000000000000000", 7383 => "0000000000000000", 7384 => "0000000000000000", 7385 => "0000000000000000", 7386 => "0000000000000000", 7387 => "0000000000000000", 7388 => "0000000000000000", 7389 => "0000000000000000", 7390 => "0000000000000000", 7391 => "0000000000000000", 7392 => "0000000000000000", 7393 => "0000000000000000", 7394 => "0000000000000000", 7395 => "0000000000000000", 7396 => "0000000000000000", 7397 => "0000000000000000", 7398 => "0000000000000000", 7399 => "0000000000000000", 7400 => "0000000000000000", 7401 => "0000000000000000", 7402 => "0000000000000000", 7403 => "0000000000000000", 7404 => "0000000000000000", 7405 => "0000000000000000", 7406 => "0000000000000000", 7407 => "0000000000000000", 7408 => "0000000000000000", 7409 => "0000000000000000", 7410 => "0000000000000000", 7411 => "0000000000000000", 7412 => "0000000000000000", 7413 => "0000000000000000", 7414 => "0000000000000000", 7415 => "0000000000000000", 7416 => "0000000000000000", 7417 => "0000000000000000", 7418 => "0000000000000000", 7419 => "0000000000000000", 7420 => "0000000000000000", 7421 => "0000000000000000", 7422 => "0000000000000000", 7423 => "0000000000000000", 7424 => "0000000000000000", 7425 => "0000000000000000", 7426 => "0000000000000000", 7427 => "0000000000000000", 7428 => "0000000000000000", 7429 => "0000000000000000", 7430 => "0000000000000000", 7431 => "0000000000000000", 7432 => "0000000000000000", 7433 => "0000000000000000", 7434 => "0000000000000000", 7435 => "0000000000000000", 7436 => "0000000000000000", 7437 => "0000000000000000", 7438 => "0000000000000000", 7439 => "0000000000000000", 7440 => "0000000000000000", 7441 => "0000000000000000", 7442 => "0000000000000000", 7443 => "0000000000000000", 7444 => "0000000000000000", 7445 => "0000000000000000", 7446 => "0000000000000000", 7447 => "0000000000000000", 7448 => "0000000000000000", 7449 => "0000000000000000", 7450 => "0000000000000000", 7451 => "0000000000000000", 7452 => "0000000000000000", 7453 => "0000000000000000", 7454 => "0000000000000000", 7455 => "0000000000000000", 7456 => "0000000000000000", 7457 => "0000000000000000", 7458 => "0000000000000000", 7459 => "0000000000000000", 7460 => "0000000000000000", 7461 => "0000000000000000", 7462 => "0000000000000000", 7463 => "0000000000000000", 7464 => "0000000000000000", 7465 => "0000000000000000", 7466 => "0000000000000000", 7467 => "0000000000000000", 7468 => "0000000000000000", 7469 => "0000000000000000", 7470 => "0000000000000000", 7471 => "0000000000000000", 7472 => "0000000000000000", 7473 => "0000000000000000", 7474 => "0000000000000000", 7475 => "0000000000000000", 7476 => "0000000000000000", 7477 => "0000000000000000", 7478 => "0000000000000000", 7479 => "0000000000000000", 7480 => "0000000000000000", 7481 => "0000000000000000", 7482 => "0000000000000000", 7483 => "0000000000000000", 7484 => "0000000000000000", 7485 => "0000000000000000", 7486 => "0000000000000000", 7487 => "0000000000000000", 7488 => "0000000000000000", 7489 => "0000000000000000", 7490 => "0000000000000000", 7491 => "0000000000000000", 7492 => "0000000000000000", 7493 => "0000000000000000", 7494 => "0000000000000000", 7495 => "0000000000000000", 7496 => "0000000000000000", 7497 => "0000000000000000", 7498 => "0000000000000000", 7499 => "0000000000000000", 7500 => "0000000000000000", 7501 => "0000000000000000", 7502 => "0000000000000000", 7503 => "0000000000000000", 7504 => "0000000000000000", 7505 => "0000000000000000", 7506 => "0000000000000000", 7507 => "0000000000000000", 7508 => "0000000000000000", 7509 => "0000000000000000", 7510 => "0000000000000000", 7511 => "0000000000000000", 7512 => "0000000000000000", 7513 => "0000000000000000", 7514 => "0000000000000000", 7515 => "0000000000000000", 7516 => "0000000000000000", 7517 => "0000000000000000", 7518 => "0000000000000000", 7519 => "0000000000000000", 7520 => "0000000000000000", 7521 => "0000000000000000", 7522 => "0000000000000000", 7523 => "0000000000000000", 7524 => "0000000000000000", 7525 => "0000000000000000", 7526 => "0000000000000000", 7527 => "0000000000000000", 7528 => "0000000000000000", 7529 => "0000000000000000", 7530 => "0000000000000000", 7531 => "0000000000000000", 7532 => "0000000000000000", 7533 => "0000000000000000", 7534 => "0000000000000000", 7535 => "0000000000000000", 7536 => "0000000000000000", 7537 => "0000000000000000", 7538 => "0000000000000000", 7539 => "0000000000000000", 7540 => "0000000000000000", 7541 => "0000000000000000", 7542 => "0000000000000000", 7543 => "0000000000000000", 7544 => "0000000000000000", 7545 => "0000000000000000", 7546 => "0000000000000000", 7547 => "0000000000000000", 7548 => "0000000000000000", 7549 => "0000000000000000", 7550 => "0000000000000000", 7551 => "0000000000000000", 7552 => "0000000000000000", 7553 => "0000000000000000", 7554 => "0000000000000000", 7555 => "0000000000000000", 7556 => "0000000000000000", 7557 => "0000000000000000", 7558 => "0000000000000000", 7559 => "0000000000000000", 7560 => "0000000000000000", 7561 => "0000000000000000", 7562 => "0000000000000000", 7563 => "0000000000000000", 7564 => "0000000000000000", 7565 => "0000000000000000", 7566 => "0000000000000000", 7567 => "0000000000000000", 7568 => "0000000000000000", 7569 => "0000000000000000", 7570 => "0000000000000000", 7571 => "0000000000000000", 7572 => "0000000000000000", 7573 => "0000000000000000", 7574 => "0000000000000000", 7575 => "0000000000000000", 7576 => "0000000000000000", 7577 => "0000000000000000", 7578 => "0000000000000000", 7579 => "0000000000000000", 7580 => "0000000000000000", 7581 => "0000000000000000", 7582 => "0000000000000000", 7583 => "0000000000000000", 7584 => "0000000000000000", 7585 => "0000000000000000", 7586 => "0000000000000000", 7587 => "0000000000000000", 7588 => "0000000000000000", 7589 => "0000000000000000", 7590 => "0000000000000000", 7591 => "0000000000000000", 7592 => "0000000000000000", 7593 => "0000000000000000", 7594 => "0000000000000000", 7595 => "0000000000000000", 7596 => "0000000000000000", 7597 => "0000000000000000", 7598 => "0000000000000000", 7599 => "0000000000000000", 7600 => "0000000000000000", 7601 => "0000000000000000", 7602 => "0000000000000000", 7603 => "0000000000000000", 7604 => "0000000000000000", 7605 => "0000000000000000", 7606 => "0000000000000000", 7607 => "0000000000000000", 7608 => "0000000000000000", 7609 => "0000000000000000", 7610 => "0000000000000000", 7611 => "0000000000000000", 7612 => "0000000000000000", 7613 => "0000000000000000", 7614 => "0000000000000000", 7615 => "0000000000000000", 7616 => "0000000000000000", 7617 => "0000000000000000", 7618 => "0000000000000000", 7619 => "0000000000000000", 7620 => "0000000000000000", 7621 => "0000000000000000", 7622 => "0000000000000000", 7623 => "0000000000000000", 7624 => "0000000000000000", 7625 => "0000000000000000", 7626 => "0000000000000000", 7627 => "0000000000000000", 7628 => "0000000000000000", 7629 => "0000000000000000", 7630 => "0000000000000000", 7631 => "0000000000000000", 7632 => "0000000000000000", 7633 => "0000000000000000", 7634 => "0000000000000000", 7635 => "0000000000000000", 7636 => "0000000000000000", 7637 => "0000000000000000", 7638 => "0000000000000000", 7639 => "0000000000000000", 7640 => "0000000000000000", 7641 => "0000000000000000", 7642 => "0000000000000000", 7643 => "0000000000000000", 7644 => "0000000000000000", 7645 => "0000000000000000", 7646 => "0000000000000000", 7647 => "0000000000000000", 7648 => "0000000000000000", 7649 => "0000000000000000", 7650 => "0000000000000000", 7651 => "0000000000000000", 7652 => "0000000000000000", 7653 => "0000000000000000", 7654 => "0000000000000000", 7655 => "0000000000000000", 7656 => "0000000000000000", 7657 => "0000000000000000", 7658 => "0000000000000000", 7659 => "0000000000000000", 7660 => "0000000000000000", 7661 => "0000000000000000", 7662 => "0000000000000000", 7663 => "0000000000000000", 7664 => "0000000000000000", 7665 => "0000000000000000", 7666 => "0000000000000000", 7667 => "0000000000000000", 7668 => "0000000000000000", 7669 => "0000000000000000", 7670 => "0000000000000000", 7671 => "0000000000000000", 7672 => "0000000000000000", 7673 => "0000000000000000", 7674 => "0000000000000000", 7675 => "0000000000000000", 7676 => "0000000000000000", 7677 => "0000000000000000", 7678 => "0000000000000000", 7679 => "0000000000000000", 7680 => "0000000000000000", 7681 => "0000000000000000", 7682 => "0000000000000000", 7683 => "0000000000000000", 7684 => "0000000000000000", 7685 => "0000000000000000", 7686 => "0000000000000000", 7687 => "0000000000000000", 7688 => "0000000000000000", 7689 => "0000000000000000", 7690 => "0000000000000000", 7691 => "0000000000000000", 7692 => "0000000000000000", 7693 => "0000000000000000", 7694 => "0000000000000000", 7695 => "0000000000000000", 7696 => "0000000000000000", 7697 => "0000000000000000", 7698 => "0000000000000000", 7699 => "0000000000000000", 7700 => "0000000000000000", 7701 => "0000000000000000", 7702 => "0000000000000000", 7703 => "0000000000000000", 7704 => "0000000000000000", 7705 => "0000000000000000", 7706 => "0000000000000000", 7707 => "0000000000000000", 7708 => "0000000000000000", 7709 => "0000000000000000", 7710 => "0000000000000000", 7711 => "0000000000000000", 7712 => "0000000000000000", 7713 => "0000000000000000", 7714 => "0000000000000000", 7715 => "0000000000000000", 7716 => "0000000000000000", 7717 => "0000000000000000", 7718 => "0000000000000000", 7719 => "0000000000000000", 7720 => "0000000000000000", 7721 => "0000000000000000", 7722 => "0000000000000000", 7723 => "0000000000000000", 7724 => "0000000000000000", 7725 => "0000000000000000", 7726 => "0000000000000000", 7727 => "0000000000000000", 7728 => "0000000000000000", 7729 => "0000000000000000", 7730 => "0000000000000000", 7731 => "0000000000000000", 7732 => "0000000000000000", 7733 => "0000000000000000", 7734 => "0000000000000000", 7735 => "0000000000000000", 7736 => "0000000000000000", 7737 => "0000000000000000", 7738 => "0000000000000000", 7739 => "0000000000000000", 7740 => "0000000000000000", 7741 => "0000000000000000", 7742 => "0000000000000000", 7743 => "0000000000000000", 7744 => "0000000000000000", 7745 => "0000000000000000", 7746 => "0000000000000000", 7747 => "0000000000000000", 7748 => "0000000000000000", 7749 => "0000000000000000", 7750 => "0000000000000000", 7751 => "0000000000000000", 7752 => "0000000000000000", 7753 => "0000000000000000", 7754 => "0000000000000000", 7755 => "0000000000000000", 7756 => "0000000000000000", 7757 => "0000000000000000", 7758 => "0000000000000000", 7759 => "0000000000000000", 7760 => "0000000000000000", 7761 => "0000000000000000", 7762 => "0000000000000000", 7763 => "0000000000000000", 7764 => "0000000000000000", 7765 => "0000000000000000", 7766 => "0000000000000000", 7767 => "0000000000000000", 7768 => "0000000000000000", 7769 => "0000000000000000", 7770 => "0000000000000000", 7771 => "0000000000000000", 7772 => "0000000000000000", 7773 => "0000000000000000", 7774 => "0000000000000000", 7775 => "0000000000000000", 7776 => "0000000000000000", 7777 => "0000000000000000", 7778 => "0000000000000000", 7779 => "0000000000000000", 7780 => "0000000000000000", 7781 => "0000000000000000", 7782 => "0000000000000000", 7783 => "0000000000000000", 7784 => "0000000000000000", 7785 => "0000000000000000", 7786 => "0000000000000000", 7787 => "0000000000000000", 7788 => "0000000000000000", 7789 => "0000000000000000", 7790 => "0000000000000000", 7791 => "0000000000000000", 7792 => "0000000000000000", 7793 => "0000000000000000", 7794 => "0000000000000000", 7795 => "0000000000000000", 7796 => "0000000000000000", 7797 => "0000000000000000", 7798 => "0000000000000000", 7799 => "0000000000000000", 7800 => "0000000000000000", 7801 => "0000000000000000", 7802 => "0000000000000000", 7803 => "0000000000000000", 7804 => "0000000000000000", 7805 => "0000000000000000", 7806 => "0000000000000000", 7807 => "0000000000000000", 7808 => "0000000000000000", 7809 => "0000000000000000", 7810 => "0000000000000000", 7811 => "0000000000000000", 7812 => "0000000000000000", 7813 => "0000000000000000", 7814 => "0000000000000000", 7815 => "0000000000000000", 7816 => "0000000000000000", 7817 => "0000000000000000", 7818 => "0000000000000000", 7819 => "0000000000000000", 7820 => "0000000000000000", 7821 => "0000000000000000", 7822 => "0000000000000000", 7823 => "0000000000000000", 7824 => "0000000000000000", 7825 => "0000000000000000", 7826 => "0000000000000000", 7827 => "0000000000000000", 7828 => "0000000000000000", 7829 => "0000000000000000", 7830 => "0000000000000000", 7831 => "0000000000000000", 7832 => "0000000000000000", 7833 => "0000000000000000", 7834 => "0000000000000000", 7835 => "0000000000000000", 7836 => "0000000000000000", 7837 => "0000000000000000", 7838 => "0000000000000000", 7839 => "0000000000000000", 7840 => "0000000000000000", 7841 => "0000000000000000", 7842 => "0000000000000000", 7843 => "0000000000000000", 7844 => "0000000000000000", 7845 => "0000000000000000", 7846 => "0000000000000000", 7847 => "0000000000000000", 7848 => "0000000000000000", 7849 => "0000000000000000", 7850 => "0000000000000000", 7851 => "0000000000000000", 7852 => "0000000000000000", 7853 => "0000000000000000", 7854 => "0000000000000000", 7855 => "0000000000000000", 7856 => "0000000000000000", 7857 => "0000000000000000", 7858 => "0000000000000000", 7859 => "0000000000000000", 7860 => "0000000000000000", 7861 => "0000000000000000", 7862 => "0000000000000000", 7863 => "0000000000000000", 7864 => "0000000000000000", 7865 => "0000000000000000", 7866 => "0000000000000000", 7867 => "0000000000000000", 7868 => "0000000000000000", 7869 => "0000000000000000", 7870 => "0000000000000000", 7871 => "0000000000000000", 7872 => "0000000000000000", 7873 => "0000000000000000", 7874 => "0000000000000000", 7875 => "0000000000000000", 7876 => "0000000000000000", 7877 => "0000000000000000", 7878 => "0000000000000000", 7879 => "0000000000000000", 7880 => "0000000000000000", 7881 => "0000000000000000", 7882 => "0000000000000000", 7883 => "0000000000000000", 7884 => "0000000000000000", 7885 => "0000000000000000", 7886 => "0000000000000000", 7887 => "0000000000000000", 7888 => "0000000000000000", 7889 => "0000000000000000", 7890 => "0000000000000000", 7891 => "0000000000000000", 7892 => "0000000000000000", 7893 => "0000000000000000", 7894 => "0000000000000000", 7895 => "0000000000000000", 7896 => "0000000000000000", 7897 => "0000000000000000", 7898 => "0000000000000000", 7899 => "0000000000000000", 7900 => "0000000000000000", 7901 => "0000000000000000", 7902 => "0000000000000000", 7903 => "0000000000000000", 7904 => "0000000000000000", 7905 => "0000000000000000", 7906 => "0000000000000000", 7907 => "0000000000000000", 7908 => "0000000000000000", 7909 => "0000000000000000", 7910 => "0000000000000000", 7911 => "0000000000000000", 7912 => "0000000000000000", 7913 => "0000000000000000", 7914 => "0000000000000000", 7915 => "0000000000000000", 7916 => "0000000000000000", 7917 => "0000000000000000", 7918 => "0000000000000000", 7919 => "0000000000000000", 7920 => "0000000000000000", 7921 => "0000000000000000", 7922 => "0000000000000000", 7923 => "0000000000000000", 7924 => "0000000000000000", 7925 => "0000000000000000", 7926 => "0000000000000000", 7927 => "0000000000000000", 7928 => "0000000000000000", 7929 => "0000000000000000", 7930 => "0000000000000000", 7931 => "0000000000000000", 7932 => "0000000000000000", 7933 => "0000000000000000", 7934 => "0000000000000000", 7935 => "0000000000000000", 7936 => "0000000000000000", 7937 => "0000000000000000", 7938 => "0000000000000000", 7939 => "0000000000000000", 7940 => "0000000000000000", 7941 => "0000000000000000", 7942 => "0000000000000000", 7943 => "0000000000000000", 7944 => "0000000000000000", 7945 => "0000000000000000", 7946 => "0000000000000000", 7947 => "0000000000000000", 7948 => "0000000000000000", 7949 => "0000000000000000", 7950 => "0000000000000000", 7951 => "0000000000000000", 7952 => "0000000000000000", 7953 => "0000000000000000", 7954 => "0000000000000000", 7955 => "0000000000000000", 7956 => "0000000000000000", 7957 => "0000000000000000", 7958 => "0000000000000000", 7959 => "0000000000000000", 7960 => "0000000000000000", 7961 => "0000000000000000", 7962 => "0000000000000000", 7963 => "0000000000000000", 7964 => "0000000000000000", 7965 => "0000000000000000", 7966 => "0000000000000000", 7967 => "0000000000000000", 7968 => "0000000000000000", 7969 => "0000000000000000", 7970 => "0000000000000000", 7971 => "0000000000000000", 7972 => "0000000000000000", 7973 => "0000000000000000", 7974 => "0000000000000000", 7975 => "0000000000000000", 7976 => "0000000000000000", 7977 => "0000000000000000", 7978 => "0000000000000000", 7979 => "0000000000000000", 7980 => "0000000000000000", 7981 => "0000000000000000", 7982 => "0000000000000000", 7983 => "0000000000000000", 7984 => "0000000000000000", 7985 => "0000000000000000", 7986 => "0000000000000000", 7987 => "0000000000000000", 7988 => "0000000000000000", 7989 => "0000000000000000", 7990 => "0000000000000000", 7991 => "0000000000000000", 7992 => "0000000000000000", 7993 => "0000000000000000", 7994 => "0000000000000000", 7995 => "0000000000000000", 7996 => "0000000000000000", 7997 => "0000000000000000", 7998 => "0000000000000000", 7999 => "0000000000000000", 8000 => "0000000000000000", 8001 => "0000000000000000", 8002 => "0000000000000000", 8003 => "0000000000000000", 8004 => "0000000000000000", 8005 => "0000000000000000", 8006 => "0000000000000000", 8007 => "0000000000000000", 8008 => "0000000000000000", 8009 => "0000000000000000", 8010 => "0000000000000000", 8011 => "0000000000000000", 8012 => "0000000000000000", 8013 => "0000000000000000", 8014 => "0000000000000000", 8015 => "0000000000000000", 8016 => "0000000000000000", 8017 => "0000000000000000", 8018 => "0000000000000000", 8019 => "0000000000000000", 8020 => "0000000000000000", 8021 => "0000000000000000", 8022 => "0000000000000000", 8023 => "0000000000000000", 8024 => "0000000000000000", 8025 => "0000000000000000", 8026 => "0000000000000000", 8027 => "0000000000000000", 8028 => "0000000000000000", 8029 => "0000000000000000", 8030 => "0000000000000000", 8031 => "0000000000000000", 8032 => "0000000000000000", 8033 => "0000000000000000", 8034 => "0000000000000000", 8035 => "0000000000000000", 8036 => "0000000000000000", 8037 => "0000000000000000", 8038 => "0000000000000000", 8039 => "0000000000000000", 8040 => "0000000000000000", 8041 => "0000000000000000", 8042 => "0000000000000000", 8043 => "0000000000000000", 8044 => "0000000000000000", 8045 => "0000000000000000", 8046 => "0000000000000000", 8047 => "0000000000000000", 8048 => "0000000000000000", 8049 => "0000000000000000", 8050 => "0000000000000000", 8051 => "0000000000000000", 8052 => "0000000000000000", 8053 => "0000000000000000", 8054 => "0000000000000000", 8055 => "0000000000000000", 8056 => "0000000000000000", 8057 => "0000000000000000", 8058 => "0000000000000000", 8059 => "0000000000000000", 8060 => "0000000000000000", 8061 => "0000000000000000", 8062 => "0000000000000000", 8063 => "0000000000000000", 8064 => "0000000000000000", 8065 => "0000000000000000", 8066 => "0000000000000000", 8067 => "0000000000000000", 8068 => "0000000000000000", 8069 => "0000000000000000", 8070 => "0000000000000000", 8071 => "0000000000000000", 8072 => "0000000000000000", 8073 => "0000000000000000", 8074 => "0000000000000000", 8075 => "0000000000000000", 8076 => "0000000000000000", 8077 => "0000000000000000", 8078 => "0000000000000000", 8079 => "0000000000000000", 8080 => "0000000000000000", 8081 => "0000000000000000", 8082 => "0000000000000000", 8083 => "0000000000000000", 8084 => "0000000000000000", 8085 => "0000000000000000", 8086 => "0000000000000000", 8087 => "0000000000000000", 8088 => "0000000000000000", 8089 => "0000000000000000", 8090 => "0000000000000000", 8091 => "0000000000000000", 8092 => "0000000000000000", 8093 => "0000000000000000", 8094 => "0000000000000000", 8095 => "0000000000000000", 8096 => "0000000000000000", 8097 => "0000000000000000", 8098 => "0000000000000000", 8099 => "0000000000000000", 8100 => "0000000000000000", 8101 => "0000000000000000", 8102 => "0000000000000000", 8103 => "0000000000000000", 8104 => "0000000000000000", 8105 => "0000000000000000", 8106 => "0000000000000000", 8107 => "0000000000000000", 8108 => "0000000000000000", 8109 => "0000000000000000", 8110 => "0000000000000000", 8111 => "0000000000000000", 8112 => "0000000000000000", 8113 => "0000000000000000", 8114 => "0000000000000000", 8115 => "0000000000000000", 8116 => "0000000000000000", 8117 => "0000000000000000", 8118 => "0000000000000000", 8119 => "0000000000000000", 8120 => "0000000000000000", 8121 => "0000000000000000", 8122 => "0000000000000000", 8123 => "0000000000000000", 8124 => "0000000000000000", 8125 => "0000000000000000", 8126 => "0000000000000000", 8127 => "0000000000000000", 8128 => "0000000000000000", 8129 => "0000000000000000", 8130 => "0000000000000000", 8131 => "0000000000000000", 8132 => "0000000000000000", 8133 => "0000000000000000", 8134 => "0000000000000000", 8135 => "0000000000000000", 8136 => "0000000000000000", 8137 => "0000000000000000", 8138 => "0000000000000000", 8139 => "0000000000000000", 8140 => "0000000000000000", 8141 => "0000000000000000", 8142 => "0000000000000000", 8143 => "0000000000000000", 8144 => "0000000000000000", 8145 => "0000000000000000", 8146 => "0000000000000000", 8147 => "0000000000000000", 8148 => "0000000000000000", 8149 => "0000000000000000", 8150 => "0000000000000000", 8151 => "0000000000000000", 8152 => "0000000000000000", 8153 => "0000000000000000", 8154 => "0000000000000000", 8155 => "0000000000000000", 8156 => "0000000000000000", 8157 => "0000000000000000", 8158 => "0000000000000000", 8159 => "0000000000000000", 8160 => "0000000000000000", 8161 => "0000000000000000", 8162 => "0000000000000000", 8163 => "0000000000000000", 8164 => "0000000000000000", 8165 => "0000000000000000", 8166 => "0000000000000000", 8167 => "0000000000000000", 8168 => "0000000000000000", 8169 => "0000000000000000", 8170 => "0000000000000000", 8171 => "0000000000000000", 8172 => "0000000000000000", 8173 => "0000000000000000", 8174 => "0000000000000000", 8175 => "0000000000000000", 8176 => "0000000000000000", 8177 => "0000000000000000", 8178 => "0000000000000000", 8179 => "0000000000000000", 8180 => "0000000000000000", 8181 => "0000000000000000", 8182 => "0000000000000000", 8183 => "0000000000000000", 8184 => "0000000000000000", 8185 => "0000000000000000", 8186 => "0000000000000000", 8187 => "0000000000000000", 8188 => "0000000000000000", 8189 => "0000000000000000", 8190 => "0000000000000000", 8191 => "0000000000000000", 8192 => "0000000000000000", 8193 => "0000000000000000", 8194 => "0000000000000000", 8195 => "0000000000000000", 8196 => "0000000000000000", 8197 => "0000000000000000", 8198 => "0000000000000000", 8199 => "0000000000000000", 8200 => "0000000000000000", 8201 => "0000000000000000", 8202 => "0000000000000000", 8203 => "0000000000000000", 8204 => "0000000000000000", 8205 => "0000000000000000", 8206 => "0000000000000000", 8207 => "0000000000000000", 8208 => "0000000000000000", 8209 => "0000000000000000", 8210 => "0000000000000000", 8211 => "0000000000000000", 8212 => "0000000000000000", 8213 => "0000000000000000", 8214 => "0000000000000000", 8215 => "0000000000000000", 8216 => "0000000000000000", 8217 => "0000000000000000", 8218 => "0000000000000000", 8219 => "0000000000000000", 8220 => "0000000000000000", 8221 => "0000000000000000", 8222 => "0000000000000000", 8223 => "0000000000000000", 8224 => "0000000000000000", 8225 => "0000000000000000", 8226 => "0000000000000000", 8227 => "0000000000000000", 8228 => "0000000000000000", 8229 => "0000000000000000", 8230 => "0000000000000000", 8231 => "0000000000000000", 8232 => "0000000000000000", 8233 => "0000000000000000", 8234 => "0000000000000000", 8235 => "0000000000000000", 8236 => "0000000000000000", 8237 => "0000000000000000", 8238 => "0000000000000000", 8239 => "0000000000000000", 8240 => "0000000000000000", 8241 => "0000000000000000", 8242 => "0000000000000000", 8243 => "0000000000000000", 8244 => "0000000000000000", 8245 => "0000000000000000", 8246 => "0000000000000000", 8247 => "0000000000000000", 8248 => "0000000000000000", 8249 => "0000000000000000", 8250 => "0000000000000000", 8251 => "0000000000000000", 8252 => "0000000000000000", 8253 => "0000000000000000", 8254 => "0000000000000000", 8255 => "0000000000000000", 8256 => "0000000000000000", 8257 => "0000000000000000", 8258 => "0000000000000000", 8259 => "0000000000000000", 8260 => "0000000000000000", 8261 => "0000000000000000", 8262 => "0000000000000000", 8263 => "0000000000000000", 8264 => "0000000000000000", 8265 => "0000000000000000", 8266 => "0000000000000000", 8267 => "0000000000000000", 8268 => "0000000000000000", 8269 => "0000000000000000", 8270 => "0000000000000000", 8271 => "0000000000000000", 8272 => "0000000000000000", 8273 => "0000000000000000", 8274 => "0000000000000000", 8275 => "0000000000000000", 8276 => "0000000000000000", 8277 => "0000000000000000", 8278 => "0000000000000000", 8279 => "0000000000000000", 8280 => "0000000000000000", 8281 => "0000000000000000", 8282 => "0000000000000000", 8283 => "0000000000000000", 8284 => "0000000000000000", 8285 => "0000000000000000", 8286 => "0000000000000000", 8287 => "0000000000000000", 8288 => "0000000000000000", 8289 => "0000000000000000", 8290 => "0000000000000000", 8291 => "0000000000000000", 8292 => "0000000000000000", 8293 => "0000000000000000", 8294 => "0000000000000000", 8295 => "0000000000000000", 8296 => "0000000000000000", 8297 => "0000000000000000", 8298 => "0000000000000000", 8299 => "0000000000000000", 8300 => "0000000000000000", 8301 => "0000000000000000", 8302 => "0000000000000000", 8303 => "0000000000000000", 8304 => "0000000000000000", 8305 => "0000000000000000", 8306 => "0000000000000000", 8307 => "0000000000000000", 8308 => "0000000000000000", 8309 => "0000000000000000", 8310 => "0000000000000000", 8311 => "0000000000000000", 8312 => "0000000000000000", 8313 => "0000000000000000", 8314 => "0000000000000000", 8315 => "0000000000000000", 8316 => "0000000000000000", 8317 => "0000000000000000", 8318 => "0000000000000000", 8319 => "0000000000000000", 8320 => "0000000000000000", 8321 => "0000000000000000", 8322 => "0000000000000000", 8323 => "0000000000000000", 8324 => "0000000000000000", 8325 => "0000000000000000", 8326 => "0000000000000000", 8327 => "0000000000000000", 8328 => "0000000000000000", 8329 => "0000000000000000", 8330 => "0000000000000000", 8331 => "0000000000000000", 8332 => "0000000000000000", 8333 => "0000000000000000", 8334 => "0000000000000000", 8335 => "0000000000000000", 8336 => "0000000000000000", 8337 => "0000000000000000", 8338 => "0000000000000000", 8339 => "0000000000000000", 8340 => "0000000000000000", 8341 => "0000000000000000", 8342 => "0000000000000000", 8343 => "0000000000000000", 8344 => "0000000000000000", 8345 => "0000000000000000", 8346 => "0000000000000000", 8347 => "0000000000000000", 8348 => "0000000000000000", 8349 => "0000000000000000", 8350 => "0000000000000000", 8351 => "0000000000000000", 8352 => "0000000000000000", 8353 => "0000000000000000", 8354 => "0000000000000000", 8355 => "0000000000000000", 8356 => "0000000000000000", 8357 => "0000000000000000", 8358 => "0000000000000000", 8359 => "0000000000000000", 8360 => "0000000000000000", 8361 => "0000000000000000", 8362 => "0000000000000000", 8363 => "0000000000000000", 8364 => "0000000000000000", 8365 => "0000000000000000", 8366 => "0000000000000000", 8367 => "0000000000000000", 8368 => "0000000000000000", 8369 => "0000000000000000", 8370 => "0000000000000000", 8371 => "0000000000000000", 8372 => "0000000000000000", 8373 => "0000000000000000", 8374 => "0000000000000000", 8375 => "0000000000000000", 8376 => "0000000000000000", 8377 => "0000000000000000", 8378 => "0000000000000000", 8379 => "0000000000000000", 8380 => "0000000000000000", 8381 => "0000000000000000", 8382 => "0000000000000000", 8383 => "0000000000000000", 8384 => "0000000000000000", 8385 => "0000000000000000", 8386 => "0000000000000000", 8387 => "0000000000000000", 8388 => "0000000000000000", 8389 => "0000000000000000", 8390 => "0000000000000000", 8391 => "0000000000000000", 8392 => "0000000000000000", 8393 => "0000000000000000", 8394 => "0000000000000000", 8395 => "0000000000000000", 8396 => "0000000000000000", 8397 => "0000000000000000", 8398 => "0000000000000000", 8399 => "0000000000000000", 8400 => "0000000000000000", 8401 => "0000000000000000", 8402 => "0000000000000000", 8403 => "0000000000000000", 8404 => "0000000000000000", 8405 => "0000000000000000", 8406 => "0000000000000000", 8407 => "0000000000000000", 8408 => "0000000000000000", 8409 => "0000000000000000", 8410 => "0000000000000000", 8411 => "0000000000000000", 8412 => "0000000000000000", 8413 => "0000000000000000", 8414 => "0000000000000000", 8415 => "0000000000000000", 8416 => "0000000000000000", 8417 => "0000000000000000", 8418 => "0000000000000000", 8419 => "0000000000000000", 8420 => "0000000000000000", 8421 => "0000000000000000", 8422 => "0000000000000000", 8423 => "0000000000000000", 8424 => "0000000000000000", 8425 => "0000000000000000", 8426 => "0000000000000000", 8427 => "0000000000000000", 8428 => "0000000000000000", 8429 => "0000000000000000", 8430 => "0000000000000000", 8431 => "0000000000000000", 8432 => "0000000000000000", 8433 => "0000000000000000", 8434 => "0000000000000000", 8435 => "0000000000000000", 8436 => "0000000000000000", 8437 => "0000000000000000", 8438 => "0000000000000000", 8439 => "0000000000000000", 8440 => "0000000000000000", 8441 => "0000000000000000", 8442 => "0000000000000000", 8443 => "0000000000000000", 8444 => "0000000000000000", 8445 => "0000000000000000", 8446 => "0000000000000000", 8447 => "0000000000000000", 8448 => "0000000000000000", 8449 => "0000000000000000", 8450 => "0000000000000000", 8451 => "0000000000000000", 8452 => "0000000000000000", 8453 => "0000000000000000", 8454 => "0000000000000000", 8455 => "0000000000000000", 8456 => "0000000000000000", 8457 => "0000000000000000", 8458 => "0000000000000000", 8459 => "0000000000000000", 8460 => "0000000000000000", 8461 => "0000000000000000", 8462 => "0000000000000000", 8463 => "0000000000000000", 8464 => "0000000000000000", 8465 => "0000000000000000", 8466 => "0000000000000000", 8467 => "0000000000000000", 8468 => "0000000000000000", 8469 => "0000000000000000", 8470 => "0000000000000000", 8471 => "0000000000000000", 8472 => "0000000000000000", 8473 => "0000000000000000", 8474 => "0000000000000000", 8475 => "0000000000000000", 8476 => "0000000000000000", 8477 => "0000000000000000", 8478 => "0000000000000000", 8479 => "0000000000000000", 8480 => "0000000000000000", 8481 => "0000000000000000", 8482 => "0000000000000000", 8483 => "0000000000000000", 8484 => "0000000000000000", 8485 => "0000000000000000", 8486 => "0000000000000000", 8487 => "0000000000000000", 8488 => "0000000000000000", 8489 => "0000000000000000", 8490 => "0000000000000000", 8491 => "0000000000000000", 8492 => "0000000000000000", 8493 => "0000000000000000", 8494 => "0000000000000000", 8495 => "0000000000000000", 8496 => "0000000000000000", 8497 => "0000000000000000", 8498 => "0000000000000000", 8499 => "0000000000000000", 8500 => "0000000000000000", 8501 => "0000000000000000", 8502 => "0000000000000000", 8503 => "0000000000000000", 8504 => "0000000000000000", 8505 => "0000000000000000", 8506 => "0000000000000000", 8507 => "0000000000000000", 8508 => "0000000000000000", 8509 => "0000000000000000", 8510 => "0000000000000000", 8511 => "0000000000000000", 8512 => "0000000000000000", 8513 => "0000000000000000", 8514 => "0000000000000000", 8515 => "0000000000000000", 8516 => "0000000000000000", 8517 => "0000000000000000", 8518 => "0000000000000000", 8519 => "0000000000000000", 8520 => "0000000000000000", 8521 => "0000000000000000", 8522 => "0000000000000000", 8523 => "0000000000000000", 8524 => "0000000000000000", 8525 => "0000000000000000", 8526 => "0000000000000000", 8527 => "0000000000000000", 8528 => "0000000000000000", 8529 => "0000000000000000", 8530 => "0000000000000000", 8531 => "0000000000000000", 8532 => "0000000000000000", 8533 => "0000000000000000", 8534 => "0000000000000000", 8535 => "0000000000000000", 8536 => "0000000000000000", 8537 => "0000000000000000", 8538 => "0000000000000000", 8539 => "0000000000000000", 8540 => "0000000000000000", 8541 => "0000000000000000", 8542 => "0000000000000000", 8543 => "0000000000000000", 8544 => "0000000000000000", 8545 => "0000000000000000", 8546 => "0000000000000000", 8547 => "0000000000000000", 8548 => "0000000000000000", 8549 => "0000000000000000", 8550 => "0000000000000000", 8551 => "0000000000000000", 8552 => "0000000000000000", 8553 => "0000000000000000", 8554 => "0000000000000000", 8555 => "0000000000000000", 8556 => "0000000000000000", 8557 => "0000000000000000", 8558 => "0000000000000000", 8559 => "0000000000000000", 8560 => "0000000000000000", 8561 => "0000000000000000", 8562 => "0000000000000000", 8563 => "0000000000000000", 8564 => "0000000000000000", 8565 => "0000000000000000", 8566 => "0000000000000000", 8567 => "0000000000000000", 8568 => "0000000000000000", 8569 => "0000000000000000", 8570 => "0000000000000000", 8571 => "0000000000000000", 8572 => "0000000000000000", 8573 => "0000000000000000", 8574 => "0000000000000000", 8575 => "0000000000000000", 8576 => "0000000000000000", 8577 => "0000000000000000", 8578 => "0000000000000000", 8579 => "0000000000000000", 8580 => "0000000000000000", 8581 => "0000000000000000", 8582 => "0000000000000000", 8583 => "0000000000000000", 8584 => "0000000000000000", 8585 => "0000000000000000", 8586 => "0000000000000000", 8587 => "0000000000000000", 8588 => "0000000000000000", 8589 => "0000000000000000", 8590 => "0000000000000000", 8591 => "0000000000000000", 8592 => "0000000000000000", 8593 => "0000000000000000", 8594 => "0000000000000000", 8595 => "0000000000000000", 8596 => "0000000000000000", 8597 => "0000000000000000", 8598 => "0000000000000000", 8599 => "0000000000000000", 8600 => "0000000000000000", 8601 => "0000000000000000", 8602 => "0000000000000000", 8603 => "0000000000000000", 8604 => "0000000000000000", 8605 => "0000000000000000", 8606 => "0000000000000000", 8607 => "0000000000000000", 8608 => "0000000000000000", 8609 => "0000000000000000", 8610 => "0000000000000000", 8611 => "0000000000000000", 8612 => "0000000000000000", 8613 => "0000000000000000", 8614 => "0000000000000000", 8615 => "0000000000000000", 8616 => "0000000000000000", 8617 => "0000000000000000", 8618 => "0000000000000000", 8619 => "0000000000000000", 8620 => "0000000000000000", 8621 => "0000000000000000", 8622 => "0000000000000000", 8623 => "0000000000000000", 8624 => "0000000000000000", 8625 => "0000000000000000", 8626 => "0000000000000000", 8627 => "0000000000000000", 8628 => "0000000000000000", 8629 => "0000000000000000", 8630 => "0000000000000000", 8631 => "0000000000000000", 8632 => "0000000000000000", 8633 => "0000000000000000", 8634 => "0000000000000000", 8635 => "0000000000000000", 8636 => "0000000000000000", 8637 => "0000000000000000", 8638 => "0000000000000000", 8639 => "0000000000000000", 8640 => "0000000000000000", 8641 => "0000000000000000", 8642 => "0000000000000000", 8643 => "0000000000000000", 8644 => "0000000000000000", 8645 => "0000000000000000", 8646 => "0000000000000000", 8647 => "0000000000000000", 8648 => "0000000000000000", 8649 => "0000000000000000", 8650 => "0000000000000000", 8651 => "0000000000000000", 8652 => "0000000000000000", 8653 => "0000000000000000", 8654 => "0000000000000000", 8655 => "0000000000000000", 8656 => "0000000000000000", 8657 => "0000000000000000", 8658 => "0000000000000000", 8659 => "0000000000000000", 8660 => "0000000000000000", 8661 => "0000000000000000", 8662 => "0000000000000000", 8663 => "0000000000000000", 8664 => "0000000000000000", 8665 => "0000000000000000", 8666 => "0000000000000000", 8667 => "0000000000000000", 8668 => "0000000000000000", 8669 => "0000000000000000", 8670 => "0000000000000000", 8671 => "0000000000000000", 8672 => "0000000000000000", 8673 => "0000000000000000", 8674 => "0000000000000000", 8675 => "0000000000000000", 8676 => "0000000000000000", 8677 => "0000000000000000", 8678 => "0000000000000000", 8679 => "0000000000000000", 8680 => "0000000000000000", 8681 => "0000000000000000", 8682 => "0000000000000000", 8683 => "0000000000000000", 8684 => "0000000000000000", 8685 => "0000000000000000", 8686 => "0000000000000000", 8687 => "0000000000000000", 8688 => "0000000000000000", 8689 => "0000000000000000", 8690 => "0000000000000000", 8691 => "0000000000000000", 8692 => "0000000000000000", 8693 => "0000000000000000", 8694 => "0000000000000000", 8695 => "0000000000000000", 8696 => "0000000000000000", 8697 => "0000000000000000", 8698 => "0000000000000000", 8699 => "0000000000000000", 8700 => "0000000000000000", 8701 => "0000000000000000", 8702 => "0000000000000000", 8703 => "0000000000000000", 8704 => "0000000000000000", 8705 => "0000000000000000", 8706 => "0000000000000000", 8707 => "0000000000000000", 8708 => "0000000000000000", 8709 => "0000000000000000", 8710 => "0000000000000000", 8711 => "0000000000000000", 8712 => "0000000000000000", 8713 => "0000000000000000", 8714 => "0000000000000000", 8715 => "0000000000000000", 8716 => "0000000000000000", 8717 => "0000000000000000", 8718 => "0000000000000000", 8719 => "0000000000000000", 8720 => "0000000000000000", 8721 => "0000000000000000", 8722 => "0000000000000000", 8723 => "0000000000000000", 8724 => "0000000000000000", 8725 => "0000000000000000", 8726 => "0000000000000000", 8727 => "0000000000000000", 8728 => "0000000000000000", 8729 => "0000000000000000", 8730 => "0000000000000000", 8731 => "0000000000000000", 8732 => "0000000000000000", 8733 => "0000000000000000", 8734 => "0000000000000000", 8735 => "0000000000000000", 8736 => "0000000000000000", 8737 => "0000000000000000", 8738 => "0000000000000000", 8739 => "0000000000000000", 8740 => "0000000000000000", 8741 => "0000000000000000", 8742 => "0000000000000000", 8743 => "0000000000000000", 8744 => "0000000000000000", 8745 => "0000000000000000", 8746 => "0000000000000000", 8747 => "0000000000000000", 8748 => "0000000000000000", 8749 => "0000000000000000", 8750 => "0000000000000000", 8751 => "0000000000000000", 8752 => "0000000000000000", 8753 => "0000000000000000", 8754 => "0000000000000000", 8755 => "0000000000000000", 8756 => "0000000000000000", 8757 => "0000000000000000", 8758 => "0000000000000000", 8759 => "0000000000000000", 8760 => "0000000000000000", 8761 => "0000000000000000", 8762 => "0000000000000000", 8763 => "0000000000000000", 8764 => "0000000000000000", 8765 => "0000000000000000", 8766 => "0000000000000000", 8767 => "0000000000000000", 8768 => "0000000000000000", 8769 => "0000000000000000", 8770 => "0000000000000000", 8771 => "0000000000000000", 8772 => "0000000000000000", 8773 => "0000000000000000", 8774 => "0000000000000000", 8775 => "0000000000000000", 8776 => "0000000000000000", 8777 => "0000000000000000", 8778 => "0000000000000000", 8779 => "0000000000000000", 8780 => "0000000000000000", 8781 => "0000000000000000", 8782 => "0000000000000000", 8783 => "0000000000000000", 8784 => "0000000000000000", 8785 => "0000000000000000", 8786 => "0000000000000000", 8787 => "0000000000000000", 8788 => "0000000000000000", 8789 => "0000000000000000", 8790 => "0000000000000000", 8791 => "0000000000000000", 8792 => "0000000000000000", 8793 => "0000000000000000", 8794 => "0000000000000000", 8795 => "0000000000000000", 8796 => "0000000000000000", 8797 => "0000000000000000", 8798 => "0000000000000000", 8799 => "0000000000000000", 8800 => "0000000000000000", 8801 => "0000000000000000", 8802 => "0000000000000000", 8803 => "0000000000000000", 8804 => "0000000000000000", 8805 => "0000000000000000", 8806 => "0000000000000000", 8807 => "0000000000000000", 8808 => "0000000000000000", 8809 => "0000000000000000", 8810 => "0000000000000000", 8811 => "0000000000000000", 8812 => "0000000000000000", 8813 => "0000000000000000", 8814 => "0000000000000000", 8815 => "0000000000000000", 8816 => "0000000000000000", 8817 => "0000000000000000", 8818 => "0000000000000000", 8819 => "0000000000000000", 8820 => "0000000000000000", 8821 => "0000000000000000", 8822 => "0000000000000000", 8823 => "0000000000000000", 8824 => "0000000000000000", 8825 => "0000000000000000", 8826 => "0000000000000000", 8827 => "0000000000000000", 8828 => "0000000000000000", 8829 => "0000000000000000", 8830 => "0000000000000000", 8831 => "0000000000000000", 8832 => "0000000000000000", 8833 => "0000000000000000", 8834 => "0000000000000000", 8835 => "0000000000000000", 8836 => "0000000000000000", 8837 => "0000000000000000", 8838 => "0000000000000000", 8839 => "0000000000000000", 8840 => "0000000000000000", 8841 => "0000000000000000", 8842 => "0000000000000000", 8843 => "0000000000000000", 8844 => "0000000000000000", 8845 => "0000000000000000", 8846 => "0000000000000000", 8847 => "0000000000000000", 8848 => "0000000000000000", 8849 => "0000000000000000", 8850 => "0000000000000000", 8851 => "0000000000000000", 8852 => "0000000000000000", 8853 => "0000000000000000", 8854 => "0000000000000000", 8855 => "0000000000000000", 8856 => "0000000000000000", 8857 => "0000000000000000", 8858 => "0000000000000000", 8859 => "0000000000000000", 8860 => "0000000000000000", 8861 => "0000000000000000", 8862 => "0000000000000000", 8863 => "0000000000000000", 8864 => "0000000000000000", 8865 => "0000000000000000", 8866 => "0000000000000000", 8867 => "0000000000000000", 8868 => "0000000000000000", 8869 => "0000000000000000", 8870 => "0000000000000000", 8871 => "0000000000000000", 8872 => "0000000000000000", 8873 => "0000000000000000", 8874 => "0000000000000000", 8875 => "0000000000000000", 8876 => "0000000000000000", 8877 => "0000000000000000", 8878 => "0000000000000000", 8879 => "0000000000000000", 8880 => "0000000000000000", 8881 => "0000000000000000", 8882 => "0000000000000000", 8883 => "0000000000000000", 8884 => "0000000000000000", 8885 => "0000000000000000", 8886 => "0000000000000000", 8887 => "0000000000000000", 8888 => "0000000000000000", 8889 => "0000000000000000", 8890 => "0000000000000000", 8891 => "0000000000000000", 8892 => "0000000000000000", 8893 => "0000000000000000", 8894 => "0000000000000000", 8895 => "0000000000000000", 8896 => "0000000000000000", 8897 => "0000000000000000", 8898 => "0000000000000000", 8899 => "0000000000000000", 8900 => "0000000000000000", 8901 => "0000000000000000", 8902 => "0000000000000000", 8903 => "0000000000000000", 8904 => "0000000000000000", 8905 => "0000000000000000", 8906 => "0000000000000000", 8907 => "0000000000000000", 8908 => "0000000000000000", 8909 => "0000000000000000", 8910 => "0000000000000000", 8911 => "0000000000000000", 8912 => "0000000000000000", 8913 => "0000000000000000", 8914 => "0000000000000000", 8915 => "0000000000000000", 8916 => "0000000000000000", 8917 => "0000000000000000", 8918 => "0000000000000000", 8919 => "0000000000000000", 8920 => "0000000000000000", 8921 => "0000000000000000", 8922 => "0000000000000000", 8923 => "0000000000000000", 8924 => "0000000000000000", 8925 => "0000000000000000", 8926 => "0000000000000000", 8927 => "0000000000000000", 8928 => "0000000000000000", 8929 => "0000000000000000", 8930 => "0000000000000000", 8931 => "0000000000000000", 8932 => "0000000000000000", 8933 => "0000000000000000", 8934 => "0000000000000000", 8935 => "0000000000000000", 8936 => "0000000000000000", 8937 => "0000000000000000", 8938 => "0000000000000000", 8939 => "0000000000000000", 8940 => "0000000000000000", 8941 => "0000000000000000", 8942 => "0000000000000000", 8943 => "0000000000000000", 8944 => "0000000000000000", 8945 => "0000000000000000", 8946 => "0000000000000000", 8947 => "0000000000000000", 8948 => "0000000000000000", 8949 => "0000000000000000", 8950 => "0000000000000000", 8951 => "0000000000000000", 8952 => "0000000000000000", 8953 => "0000000000000000", 8954 => "0000000000000000", 8955 => "0000000000000000", 8956 => "0000000000000000", 8957 => "0000000000000000", 8958 => "0000000000000000", 8959 => "0000000000000000", 8960 => "0000000000000000", 8961 => "0000000000000000", 8962 => "0000000000000000", 8963 => "0000000000000000", 8964 => "0000000000000000", 8965 => "0000000000000000", 8966 => "0000000000000000", 8967 => "0000000000000000", 8968 => "0000000000000000", 8969 => "0000000000000000", 8970 => "0000000000000000", 8971 => "0000000000000000", 8972 => "0000000000000000", 8973 => "0000000000000000", 8974 => "0000000000000000", 8975 => "0000000000000000", 8976 => "0000000000000000", 8977 => "0000000000000000", 8978 => "0000000000000000", 8979 => "0000000000000000", 8980 => "0000000000000000", 8981 => "0000000000000000", 8982 => "0000000000000000", 8983 => "0000000000000000", 8984 => "0000000000000000", 8985 => "0000000000000000", 8986 => "0000000000000000", 8987 => "0000000000000000", 8988 => "0000000000000000", 8989 => "0000000000000000", 8990 => "0000000000000000", 8991 => "0000000000000000", 8992 => "0000000000000000", 8993 => "0000000000000000", 8994 => "0000000000000000", 8995 => "0000000000000000", 8996 => "0000000000000000", 8997 => "0000000000000000", 8998 => "0000000000000000", 8999 => "0000000000000000", 9000 => "0000000000000000", 9001 => "0000000000000000", 9002 => "0000000000000000", 9003 => "0000000000000000", 9004 => "0000000000000000", 9005 => "0000000000000000", 9006 => "0000000000000000", 9007 => "0000000000000000", 9008 => "0000000000000000", 9009 => "0000000000000000", 9010 => "0000000000000000", 9011 => "0000000000000000", 9012 => "0000000000000000", 9013 => "0000000000000000", 9014 => "0000000000000000", 9015 => "0000000000000000", 9016 => "0000000000000000", 9017 => "0000000000000000", 9018 => "0000000000000000", 9019 => "0000000000000000", 9020 => "0000000000000000", 9021 => "0000000000000000", 9022 => "0000000000000000", 9023 => "0000000000000000", 9024 => "0000000000000000", 9025 => "0000000000000000", 9026 => "0000000000000000", 9027 => "0000000000000000", 9028 => "0000000000000000", 9029 => "0000000000000000", 9030 => "0000000000000000", 9031 => "0000000000000000", 9032 => "0000000000000000", 9033 => "0000000000000000", 9034 => "0000000000000000", 9035 => "0000000000000000", 9036 => "0000000000000000", 9037 => "0000000000000000", 9038 => "0000000000000000", 9039 => "0000000000000000", 9040 => "0000000000000000", 9041 => "0000000000000000", 9042 => "0000000000000000", 9043 => "0000000000000000", 9044 => "0000000000000000", 9045 => "0000000000000000", 9046 => "0000000000000000", 9047 => "0000000000000000", 9048 => "0000000000000000", 9049 => "0000000000000000", 9050 => "0000000000000000", 9051 => "0000000000000000", 9052 => "0000000000000000", 9053 => "0000000000000000", 9054 => "0000000000000000", 9055 => "0000000000000000", 9056 => "0000000000000000", 9057 => "0000000000000000", 9058 => "0000000000000000", 9059 => "0000000000000000", 9060 => "0000000000000000", 9061 => "0000000000000000", 9062 => "0000000000000000", 9063 => "0000000000000000", 9064 => "0000000000000000", 9065 => "0000000000000000", 9066 => "0000000000000000", 9067 => "0000000000000000", 9068 => "0000000000000000", 9069 => "0000000000000000", 9070 => "0000000000000000", 9071 => "0000000000000000", 9072 => "0000000000000000", 9073 => "0000000000000000", 9074 => "0000000000000000", 9075 => "0000000000000000", 9076 => "0000000000000000", 9077 => "0000000000000000", 9078 => "0000000000000000", 9079 => "0000000000000000", 9080 => "0000000000000000", 9081 => "0000000000000000", 9082 => "0000000000000000", 9083 => "0000000000000000", 9084 => "0000000000000000", 9085 => "0000000000000000", 9086 => "0000000000000000", 9087 => "0000000000000000", 9088 => "0000000000000000", 9089 => "0000000000000000", 9090 => "0000000000000000", 9091 => "0000000000000000", 9092 => "0000000000000000", 9093 => "0000000000000000", 9094 => "0000000000000000", 9095 => "0000000000000000", 9096 => "0000000000000000", 9097 => "0000000000000000", 9098 => "0000000000000000", 9099 => "0000000000000000", 9100 => "0000000000000000", 9101 => "0000000000000000", 9102 => "0000000000000000", 9103 => "0000000000000000", 9104 => "0000000000000000", 9105 => "0000000000000000", 9106 => "0000000000000000", 9107 => "0000000000000000", 9108 => "0000000000000000", 9109 => "0000000000000000", 9110 => "0000000000000000", 9111 => "0000000000000000", 9112 => "0000000000000000", 9113 => "0000000000000000", 9114 => "0000000000000000", 9115 => "0000000000000000", 9116 => "0000000000000000", 9117 => "0000000000000000", 9118 => "0000000000000000", 9119 => "0000000000000000", 9120 => "0000000000000000", 9121 => "0000000000000000", 9122 => "0000000000000000", 9123 => "0000000000000000", 9124 => "0000000000000000", 9125 => "0000000000000000", 9126 => "0000000000000000", 9127 => "0000000000000000", 9128 => "0000000000000000", 9129 => "0000000000000000", 9130 => "0000000000000000", 9131 => "0000000000000000", 9132 => "0000000000000000", 9133 => "0000000000000000", 9134 => "0000000000000000", 9135 => "0000000000000000", 9136 => "0000000000000000", 9137 => "0000000000000000", 9138 => "0000000000000000", 9139 => "0000000000000000", 9140 => "0000000000000000", 9141 => "0000000000000000", 9142 => "0000000000000000", 9143 => "0000000000000000", 9144 => "0000000000000000", 9145 => "0000000000000000", 9146 => "0000000000000000", 9147 => "0000000000000000", 9148 => "0000000000000000", 9149 => "0000000000000000", 9150 => "0000000000000000", 9151 => "0000000000000000", 9152 => "0000000000000000", 9153 => "0000000000000000", 9154 => "0000000000000000", 9155 => "0000000000000000", 9156 => "0000000000000000", 9157 => "0000000000000000", 9158 => "0000000000000000", 9159 => "0000000000000000", 9160 => "0000000000000000", 9161 => "0000000000000000", 9162 => "0000000000000000", 9163 => "0000000000000000", 9164 => "0000000000000000", 9165 => "0000000000000000", 9166 => "0000000000000000", 9167 => "0000000000000000", 9168 => "0000000000000000", 9169 => "0000000000000000", 9170 => "0000000000000000", 9171 => "0000000000000000", 9172 => "0000000000000000", 9173 => "0000000000000000", 9174 => "0000000000000000", 9175 => "0000000000000000", 9176 => "0000000000000000", 9177 => "0000000000000000", 9178 => "0000000000000000", 9179 => "0000000000000000", 9180 => "0000000000000000", 9181 => "0000000000000000", 9182 => "0000000000000000", 9183 => "0000000000000000", 9184 => "0000000000000000", 9185 => "0000000000000000", 9186 => "0000000000000000", 9187 => "0000000000000000", 9188 => "0000000000000000", 9189 => "0000000000000000", 9190 => "0000000000000000", 9191 => "0000000000000000", 9192 => "0000000000000000", 9193 => "0000000000000000", 9194 => "0000000000000000", 9195 => "0000000000000000", 9196 => "0000000000000000", 9197 => "0000000000000000", 9198 => "0000000000000000", 9199 => "0000000000000000", 9200 => "0000000000000000", 9201 => "0000000000000000", 9202 => "0000000000000000", 9203 => "0000000000000000", 9204 => "0000000000000000", 9205 => "0000000000000000", 9206 => "0000000000000000", 9207 => "0000000000000000", 9208 => "0000000000000000", 9209 => "0000000000000000", 9210 => "0000000000000000", 9211 => "0000000000000000", 9212 => "0000000000000000", 9213 => "0000000000000000", 9214 => "0000000000000000", 9215 => "0000000000000000", 9216 => "0000000000000000", 9217 => "0000000000000000", 9218 => "0000000000000000", 9219 => "0000000000000000", 9220 => "0000000000000000", 9221 => "0000000000000000", 9222 => "0000000000000000", 9223 => "0000000000000000", 9224 => "0000000000000000", 9225 => "0000000000000000", 9226 => "0000000000000000", 9227 => "0000000000000000", 9228 => "0000000000000000", 9229 => "0000000000000000", 9230 => "0000000000000000", 9231 => "0000000000000000", 9232 => "0000000000000000", 9233 => "0000000000000000", 9234 => "0000000000000000", 9235 => "0000000000000000", 9236 => "0000000000000000", 9237 => "0000000000000000", 9238 => "0000000000000000", 9239 => "0000000000000000", 9240 => "0000000000000000", 9241 => "0000000000000000", 9242 => "0000000000000000", 9243 => "0000000000000000", 9244 => "0000000000000000", 9245 => "0000000000000000", 9246 => "0000000000000000", 9247 => "0000000000000000", 9248 => "0000000000000000", 9249 => "0000000000000000", 9250 => "0000000000000000", 9251 => "0000000000000000", 9252 => "0000000000000000", 9253 => "0000000000000000", 9254 => "0000000000000000", 9255 => "0000000000000000", 9256 => "0000000000000000", 9257 => "0000000000000000", 9258 => "0000000000000000", 9259 => "0000000000000000", 9260 => "0000000000000000", 9261 => "0000000000000000", 9262 => "0000000000000000", 9263 => "0000000000000000", 9264 => "0000000000000000", 9265 => "0000000000000000", 9266 => "0000000000000000", 9267 => "0000000000000000", 9268 => "0000000000000000", 9269 => "0000000000000000", 9270 => "0000000000000000", 9271 => "0000000000000000", 9272 => "0000000000000000", 9273 => "0000000000000000", 9274 => "0000000000000000", 9275 => "0000000000000000", 9276 => "0000000000000000", 9277 => "0000000000000000", 9278 => "0000000000000000", 9279 => "0000000000000000", 9280 => "0000000000000000", 9281 => "0000000000000000", 9282 => "0000000000000000", 9283 => "0000000000000000", 9284 => "0000000000000000", 9285 => "0000000000000000", 9286 => "0000000000000000", 9287 => "0000000000000000", 9288 => "0000000000000000", 9289 => "0000000000000000", 9290 => "0000000000000000", 9291 => "0000000000000000", 9292 => "0000000000000000", 9293 => "0000000000000000", 9294 => "0000000000000000", 9295 => "0000000000000000", 9296 => "0000000000000000", 9297 => "0000000000000000", 9298 => "0000000000000000", 9299 => "0000000000000000", 9300 => "0000000000000000", 9301 => "0000000000000000", 9302 => "0000000000000000", 9303 => "0000000000000000", 9304 => "0000000000000000", 9305 => "0000000000000000", 9306 => "0000000000000000", 9307 => "0000000000000000", 9308 => "0000000000000000", 9309 => "0000000000000000", 9310 => "0000000000000000", 9311 => "0000000000000000", 9312 => "0000000000000000", 9313 => "0000000000000000", 9314 => "0000000000000000", 9315 => "0000000000000000", 9316 => "0000000000000000", 9317 => "0000000000000000", 9318 => "0000000000000000", 9319 => "0000000000000000", 9320 => "0000000000000000", 9321 => "0000000000000000", 9322 => "0000000000000000", 9323 => "0000000000000000", 9324 => "0000000000000000", 9325 => "0000000000000000", 9326 => "0000000000000000", 9327 => "0000000000000000", 9328 => "0000000000000000", 9329 => "0000000000000000", 9330 => "0000000000000000", 9331 => "0000000000000000", 9332 => "0000000000000000", 9333 => "0000000000000000", 9334 => "0000000000000000", 9335 => "0000000000000000", 9336 => "0000000000000000", 9337 => "0000000000000000", 9338 => "0000000000000000", 9339 => "0000000000000000", 9340 => "0000000000000000", 9341 => "0000000000000000", 9342 => "0000000000000000", 9343 => "0000000000000000", 9344 => "0000000000000000", 9345 => "0000000000000000", 9346 => "0000000000000000", 9347 => "0000000000000000", 9348 => "0000000000000000", 9349 => "0000000000000000", 9350 => "0000000000000000", 9351 => "0000000000000000", 9352 => "0000000000000000", 9353 => "0000000000000000", 9354 => "0000000000000000", 9355 => "0000000000000000", 9356 => "0000000000000000", 9357 => "0000000000000000", 9358 => "0000000000000000", 9359 => "0000000000000000", 9360 => "0000000000000000", 9361 => "0000000000000000", 9362 => "0000000000000000", 9363 => "0000000000000000", 9364 => "0000000000000000", 9365 => "0000000000000000", 9366 => "0000000000000000", 9367 => "0000000000000000", 9368 => "0000000000000000", 9369 => "0000000000000000", 9370 => "0000000000000000", 9371 => "0000000000000000", 9372 => "0000000000000000", 9373 => "0000000000000000", 9374 => "0000000000000000", 9375 => "0000000000000000", 9376 => "0000000000000000", 9377 => "0000000000000000", 9378 => "0000000000000000", 9379 => "0000000000000000", 9380 => "0000000000000000", 9381 => "0000000000000000", 9382 => "0000000000000000", 9383 => "0000000000000000", 9384 => "0000000000000000", 9385 => "0000000000000000", 9386 => "0000000000000000", 9387 => "0000000000000000", 9388 => "0000000000000000", 9389 => "0000000000000000", 9390 => "0000000000000000", 9391 => "0000000000000000", 9392 => "0000000000000000", 9393 => "0000000000000000", 9394 => "0000000000000000", 9395 => "0000000000000000", 9396 => "0000000000000000", 9397 => "0000000000000000", 9398 => "0000000000000000", 9399 => "0000000000000000", 9400 => "0000000000000000", 9401 => "0000000000000000", 9402 => "0000000000000000", 9403 => "0000000000000000", 9404 => "0000000000000000", 9405 => "0000000000000000", 9406 => "0000000000000000", 9407 => "0000000000000000", 9408 => "0000000000000000", 9409 => "0000000000000000", 9410 => "0000000000000000", 9411 => "0000000000000000", 9412 => "0000000000000000", 9413 => "0000000000000000", 9414 => "0000000000000000", 9415 => "0000000000000000", 9416 => "0000000000000000", 9417 => "0000000000000000", 9418 => "0000000000000000", 9419 => "0000000000000000", 9420 => "0000000000000000", 9421 => "0000000000000000", 9422 => "0000000000000000", 9423 => "0000000000000000", 9424 => "0000000000000000", 9425 => "0000000000000000", 9426 => "0000000000000000", 9427 => "0000000000000000", 9428 => "0000000000000000", 9429 => "0000000000000000", 9430 => "0000000000000000", 9431 => "0000000000000000", 9432 => "0000000000000000", 9433 => "0000000000000000", 9434 => "0000000000000000", 9435 => "0000000000000000", 9436 => "0000000000000000", 9437 => "0000000000000000", 9438 => "0000000000000000", 9439 => "0000000000000000", 9440 => "0000000000000000", 9441 => "0000000000000000", 9442 => "0000000000000000", 9443 => "0000000000000000", 9444 => "0000000000000000", 9445 => "0000000000000000", 9446 => "0000000000000000", 9447 => "0000000000000000", 9448 => "0000000000000000", 9449 => "0000000000000000", 9450 => "0000000000000000", 9451 => "0000000000000000", 9452 => "0000000000000000", 9453 => "0000000000000000", 9454 => "0000000000000000", 9455 => "0000000000000000", 9456 => "0000000000000000", 9457 => "0000000000000000", 9458 => "0000000000000000", 9459 => "0000000000000000", 9460 => "0000000000000000", 9461 => "0000000000000000", 9462 => "0000000000000000", 9463 => "0000000000000000", 9464 => "0000000000000000", 9465 => "0000000000000000", 9466 => "0000000000000000", 9467 => "0000000000000000", 9468 => "0000000000000000", 9469 => "0000000000000000", 9470 => "0000000000000000", 9471 => "0000000000000000", 9472 => "0000000000000000", 9473 => "0000000000000000", 9474 => "0000000000000000", 9475 => "0000000000000000", 9476 => "0000000000000000", 9477 => "0000000000000000", 9478 => "0000000000000000", 9479 => "0000000000000000", 9480 => "0000000000000000", 9481 => "0000000000000000", 9482 => "0000000000000000", 9483 => "0000000000000000", 9484 => "0000000000000000", 9485 => "0000000000000000", 9486 => "0000000000000000", 9487 => "0000000000000000", 9488 => "0000000000000000", 9489 => "0000000000000000", 9490 => "0000000000000000", 9491 => "0000000000000000", 9492 => "0000000000000000", 9493 => "0000000000000000", 9494 => "0000000000000000", 9495 => "0000000000000000", 9496 => "0000000000000000", 9497 => "0000000000000000", 9498 => "0000000000000000", 9499 => "0000000000000000", 9500 => "0000000000000000", 9501 => "0000000000000000", 9502 => "0000000000000000", 9503 => "0000000000000000", 9504 => "0000000000000000", 9505 => "0000000000000000", 9506 => "0000000000000000", 9507 => "0000000000000000", 9508 => "0000000000000000", 9509 => "0000000000000000", 9510 => "0000000000000000", 9511 => "0000000000000000", 9512 => "0000000000000000", 9513 => "0000000000000000", 9514 => "0000000000000000", 9515 => "0000000000000000", 9516 => "0000000000000000", 9517 => "0000000000000000", 9518 => "0000000000000000", 9519 => "0000000000000000", 9520 => "0000000000000000", 9521 => "0000000000000000", 9522 => "0000000000000000", 9523 => "0000000000000000", 9524 => "0000000000000000", 9525 => "0000000000000000", 9526 => "0000000000000000", 9527 => "0000000000000000", 9528 => "0000000000000000", 9529 => "0000000000000000", 9530 => "0000000000000000", 9531 => "0000000000000000", 9532 => "0000000000000000", 9533 => "0000000000000000", 9534 => "0000000000000000", 9535 => "0000000000000000", 9536 => "0000000000000000", 9537 => "0000000000000000", 9538 => "0000000000000000", 9539 => "0000000000000000", 9540 => "0000000000000000", 9541 => "0000000000000000", 9542 => "0000000000000000", 9543 => "0000000000000000", 9544 => "0000000000000000", 9545 => "0000000000000000", 9546 => "0000000000000000", 9547 => "0000000000000000", 9548 => "0000000000000000", 9549 => "0000000000000000", 9550 => "0000000000000000", 9551 => "0000000000000000", 9552 => "0000000000000000", 9553 => "0000000000000000", 9554 => "0000000000000000", 9555 => "0000000000000000", 9556 => "0000000000000000", 9557 => "0000000000000000", 9558 => "0000000000000000", 9559 => "0000000000000000", 9560 => "0000000000000000", 9561 => "0000000000000000", 9562 => "0000000000000000", 9563 => "0000000000000000", 9564 => "0000000000000000", 9565 => "0000000000000000", 9566 => "0000000000000000", 9567 => "0000000000000000", 9568 => "0000000000000000", 9569 => "0000000000000000", 9570 => "0000000000000000", 9571 => "0000000000000000", 9572 => "0000000000000000", 9573 => "0000000000000000", 9574 => "0000000000000000", 9575 => "0000000000000000", 9576 => "0000000000000000", 9577 => "0000000000000000", 9578 => "0000000000000000", 9579 => "0000000000000000", 9580 => "0000000000000000", 9581 => "0000000000000000", 9582 => "0000000000000000", 9583 => "0000000000000000", 9584 => "0000000000000000", 9585 => "0000000000000000", 9586 => "0000000000000000", 9587 => "0000000000000000", 9588 => "0000000000000000", 9589 => "0000000000000000", 9590 => "0000000000000000", 9591 => "0000000000000000", 9592 => "0000000000000000", 9593 => "0000000000000000", 9594 => "0000000000000000", 9595 => "0000000000000000", 9596 => "0000000000000000", 9597 => "0000000000000000", 9598 => "0000000000000000", 9599 => "0000000000000000", 9600 => "0000000000000000", 9601 => "0000000000000000", 9602 => "0000000000000000", 9603 => "0000000000000000", 9604 => "0000000000000000", 9605 => "0000000000000000", 9606 => "0000000000000000", 9607 => "0000000000000000", 9608 => "0000000000000000", 9609 => "0000000000000000", 9610 => "0000000000000000", 9611 => "0000000000000000", 9612 => "0000000000000000", 9613 => "0000000000000000", 9614 => "0000000000000000", 9615 => "0000000000000000", 9616 => "0000000000000000", 9617 => "0000000000000000", 9618 => "0000000000000000", 9619 => "0000000000000000", 9620 => "0000000000000000", 9621 => "0000000000000000", 9622 => "0000000000000000", 9623 => "0000000000000000", 9624 => "0000000000000000", 9625 => "0000000000000000", 9626 => "0000000000000000", 9627 => "0000000000000000", 9628 => "0000000000000000", 9629 => "0000000000000000", 9630 => "0000000000000000", 9631 => "0000000000000000", 9632 => "0000000000000000", 9633 => "0000000000000000", 9634 => "0000000000000000", 9635 => "0000000000000000", 9636 => "0000000000000000", 9637 => "0000000000000000", 9638 => "0000000000000000", 9639 => "0000000000000000", 9640 => "0000000000000000", 9641 => "0000000000000000", 9642 => "0000000000000000", 9643 => "0000000000000000", 9644 => "0000000000000000", 9645 => "0000000000000000", 9646 => "0000000000000000", 9647 => "0000000000000000", 9648 => "0000000000000000", 9649 => "0000000000000000", 9650 => "0000000000000000", 9651 => "0000000000000000", 9652 => "0000000000000000", 9653 => "0000000000000000", 9654 => "0000000000000000", 9655 => "0000000000000000", 9656 => "0000000000000000", 9657 => "0000000000000000", 9658 => "0000000000000000", 9659 => "0000000000000000", 9660 => "0000000000000000", 9661 => "0000000000000000", 9662 => "0000000000000000", 9663 => "0000000000000000", 9664 => "0000000000000000", 9665 => "0000000000000000", 9666 => "0000000000000000", 9667 => "0000000000000000", 9668 => "0000000000000000", 9669 => "0000000000000000", 9670 => "0000000000000000", 9671 => "0000000000000000", 9672 => "0000000000000000", 9673 => "0000000000000000", 9674 => "0000000000000000", 9675 => "0000000000000000", 9676 => "0000000000000000", 9677 => "0000000000000000", 9678 => "0000000000000000", 9679 => "0000000000000000", 9680 => "0000000000000000", 9681 => "0000000000000000", 9682 => "0000000000000000", 9683 => "0000000000000000", 9684 => "0000000000000000", 9685 => "0000000000000000", 9686 => "0000000000000000", 9687 => "0000000000000000", 9688 => "0000000000000000", 9689 => "0000000000000000", 9690 => "0000000000000000", 9691 => "0000000000000000", 9692 => "0000000000000000", 9693 => "0000000000000000", 9694 => "0000000000000000", 9695 => "0000000000000000", 9696 => "0000000000000000", 9697 => "0000000000000000", 9698 => "0000000000000000", 9699 => "0000000000000000", 9700 => "0000000000000000", 9701 => "0000000000000000", 9702 => "0000000000000000", 9703 => "0000000000000000", 9704 => "0000000000000000", 9705 => "0000000000000000", 9706 => "0000000000000000", 9707 => "0000000000000000", 9708 => "0000000000000000", 9709 => "0000000000000000", 9710 => "0000000000000000", 9711 => "0000000000000000", 9712 => "0000000000000000", 9713 => "0000000000000000", 9714 => "0000000000000000", 9715 => "0000000000000000", 9716 => "0000000000000000", 9717 => "0000000000000000", 9718 => "0000000000000000", 9719 => "0000000000000000", 9720 => "0000000000000000", 9721 => "0000000000000000", 9722 => "0000000000000000", 9723 => "0000000000000000", 9724 => "0000000000000000", 9725 => "0000000000000000", 9726 => "0000000000000000", 9727 => "0000000000000000", 9728 => "0000000000000000", 9729 => "0000000000000000", 9730 => "0000000000000000", 9731 => "0000000000000000", 9732 => "0000000000000000", 9733 => "0000000000000000", 9734 => "0000000000000000", 9735 => "0000000000000000", 9736 => "0000000000000000", 9737 => "0000000000000000", 9738 => "0000000000000000", 9739 => "0000000000000000", 9740 => "0000000000000000", 9741 => "0000000000000000", 9742 => "0000000000000000", 9743 => "0000000000000000", 9744 => "0000000000000000", 9745 => "0000000000000000", 9746 => "0000000000000000", 9747 => "0000000000000000", 9748 => "0000000000000000", 9749 => "0000000000000000", 9750 => "0000000000000000", 9751 => "0000000000000000", 9752 => "0000000000000000", 9753 => "0000000000000000", 9754 => "0000000000000000", 9755 => "0000000000000000", 9756 => "0000000000000000", 9757 => "0000000000000000", 9758 => "0000000000000000", 9759 => "0000000000000000", 9760 => "0000000000000000", 9761 => "0000000000000000", 9762 => "0000000000000000", 9763 => "0000000000000000", 9764 => "0000000000000000", 9765 => "0000000000000000", 9766 => "0000000000000000", 9767 => "0000000000000000", 9768 => "0000000000000000", 9769 => "0000000000000000", 9770 => "0000000000000000", 9771 => "0000000000000000", 9772 => "0000000000000000", 9773 => "0000000000000000", 9774 => "0000000000000000", 9775 => "0000000000000000", 9776 => "0000000000000000", 9777 => "0000000000000000", 9778 => "0000000000000000", 9779 => "0000000000000000", 9780 => "0000000000000000", 9781 => "0000000000000000", 9782 => "0000000000000000", 9783 => "0000000000000000", 9784 => "0000000000000000", 9785 => "0000000000000000", 9786 => "0000000000000000", 9787 => "0000000000000000", 9788 => "0000000000000000", 9789 => "0000000000000000", 9790 => "0000000000000000", 9791 => "0000000000000000", 9792 => "0000000000000000", 9793 => "0000000000000000", 9794 => "0000000000000000", 9795 => "0000000000000000", 9796 => "0000000000000000", 9797 => "0000000000000000", 9798 => "0000000000000000", 9799 => "0000000000000000", 9800 => "0000000000000000", 9801 => "0000000000000000", 9802 => "0000000000000000", 9803 => "0000000000000000", 9804 => "0000000000000000", 9805 => "0000000000000000", 9806 => "0000000000000000", 9807 => "0000000000000000", 9808 => "0000000000000000", 9809 => "0000000000000000", 9810 => "0000000000000000", 9811 => "0000000000000000", 9812 => "0000000000000000", 9813 => "0000000000000000", 9814 => "0000000000000000", 9815 => "0000000000000000", 9816 => "0000000000000000", 9817 => "0000000000000000", 9818 => "0000000000000000", 9819 => "0000000000000000", 9820 => "0000000000000000", 9821 => "0000000000000000", 9822 => "0000000000000000", 9823 => "0000000000000000", 9824 => "0000000000000000", 9825 => "0000000000000000", 9826 => "0000000000000000", 9827 => "0000000000000000", 9828 => "0000000000000000", 9829 => "0000000000000000", 9830 => "0000000000000000", 9831 => "0000000000000000", 9832 => "0000000000000000", 9833 => "0000000000000000", 9834 => "0000000000000000", 9835 => "0000000000000000", 9836 => "0000000000000000", 9837 => "0000000000000000", 9838 => "0000000000000000", 9839 => "0000000000000000", 9840 => "0000000000000000", 9841 => "0000000000000000", 9842 => "0000000000000000", 9843 => "0000000000000000", 9844 => "0000000000000000", 9845 => "0000000000000000", 9846 => "0000000000000000", 9847 => "0000000000000000", 9848 => "0000000000000000", 9849 => "0000000000000000", 9850 => "0000000000000000", 9851 => "0000000000000000", 9852 => "0000000000000000", 9853 => "0000000000000000", 9854 => "0000000000000000", 9855 => "0000000000000000", 9856 => "0000000000000000", 9857 => "0000000000000000", 9858 => "0000000000000000", 9859 => "0000000000000000", 9860 => "0000000000000000", 9861 => "0000000000000000", 9862 => "0000000000000000", 9863 => "0000000000000000", 9864 => "0000000000000000", 9865 => "0000000000000000", 9866 => "0000000000000000", 9867 => "0000000000000000", 9868 => "0000000000000000", 9869 => "0000000000000000", 9870 => "0000000000000000", 9871 => "0000000000000000", 9872 => "0000000000000000", 9873 => "0000000000000000", 9874 => "0000000000000000", 9875 => "0000000000000000", 9876 => "0000000000000000", 9877 => "0000000000000000", 9878 => "0000000000000000", 9879 => "0000000000000000", 9880 => "0000000000000000", 9881 => "0000000000000000", 9882 => "0000000000000000", 9883 => "0000000000000000", 9884 => "0000000000000000", 9885 => "0000000000000000", 9886 => "0000000000000000", 9887 => "0000000000000000", 9888 => "0000000000000000", 9889 => "0000000000000000", 9890 => "0000000000000000", 9891 => "0000000000000000", 9892 => "0000000000000000", 9893 => "0000000000000000", 9894 => "0000000000000000", 9895 => "0000000000000000", 9896 => "0000000000000000", 9897 => "0000000000000000", 9898 => "0000000000000000", 9899 => "0000000000000000", 9900 => "0000000000000000", 9901 => "0000000000000000", 9902 => "0000000000000000", 9903 => "0000000000000000", 9904 => "0000000000000000", 9905 => "0000000000000000", 9906 => "0000000000000000", 9907 => "0000000000000000", 9908 => "0000000000000000", 9909 => "0000000000000000", 9910 => "0000000000000000", 9911 => "0000000000000000", 9912 => "0000000000000000", 9913 => "0000000000000000", 9914 => "0000000000000000", 9915 => "0000000000000000", 9916 => "0000000000000000", 9917 => "0000000000000000", 9918 => "0000000000000000", 9919 => "0000000000000000", 9920 => "0000000000000000", 9921 => "0000000000000000", 9922 => "0000000000000000", 9923 => "0000000000000000", 9924 => "0000000000000000", 9925 => "0000000000000000", 9926 => "0000000000000000", 9927 => "0000000000000000", 9928 => "0000000000000000", 9929 => "0000000000000000", 9930 => "0000000000000000", 9931 => "0000000000000000", 9932 => "0000000000000000", 9933 => "0000000000000000", 9934 => "0000000000000000", 9935 => "0000000000000000", 9936 => "0000000000000000", 9937 => "0000000000000000", 9938 => "0000000000000000", 9939 => "0000000000000000", 9940 => "0000000000000000", 9941 => "0000000000000000", 9942 => "0000000000000000", 9943 => "0000000000000000", 9944 => "0000000000000000", 9945 => "0000000000000000", 9946 => "0000000000000000", 9947 => "0000000000000000", 9948 => "0000000000000000", 9949 => "0000000000000000", 9950 => "0000000000000000", 9951 => "0000000000000000", 9952 => "0000000000000000", 9953 => "0000000000000000", 9954 => "0000000000000000", 9955 => "0000000000000000", 9956 => "0000000000000000", 9957 => "0000000000000000", 9958 => "0000000000000000", 9959 => "0000000000000000", 9960 => "0000000000000000", 9961 => "0000000000000000", 9962 => "0000000000000000", 9963 => "0000000000000000", 9964 => "0000000000000000", 9965 => "0000000000000000", 9966 => "0000000000000000", 9967 => "0000000000000000", 9968 => "0000000000000000", 9969 => "0000000000000000", 9970 => "0000000000000000", 9971 => "0000000000000000", 9972 => "0000000000000000", 9973 => "0000000000000000", 9974 => "0000000000000000", 9975 => "0000000000000000", 9976 => "0000000000000000", 9977 => "0000000000000000", 9978 => "0000000000000000", 9979 => "0000000000000000", 9980 => "0000000000000000", 9981 => "0000000000000000", 9982 => "0000000000000000", 9983 => "0000000000000000", 9984 => "0000000000000000", 9985 => "0000000000000000", 9986 => "0000000000000000", 9987 => "0000000000000000", 9988 => "0000000000000000", 9989 => "0000000000000000", 9990 => "0000000000000000", 9991 => "0000000000000000", 9992 => "0000000000000000", 9993 => "0000000000000000", 9994 => "0000000000000000", 9995 => "0000000000000000", 9996 => "0000000000000000", 9997 => "0000000000000000", 9998 => "0000000000000000", 9999 => "0000000000000000", 10000 => "0000000000000000", 10001 => "0000000000000000", 10002 => "0000000000000000", 10003 => "0000000000000000", 10004 => "0000000000000000", 10005 => "0000000000000000", 10006 => "0000000000000000", 10007 => "0000000000000000", 10008 => "0000000000000000", 10009 => "0000000000000000", 10010 => "0000000000000000", 10011 => "0000000000000000", 10012 => "0000000000000000", 10013 => "0000000000000000", 10014 => "0000000000000000", 10015 => "0000000000000000", 10016 => "0000000000000000", 10017 => "0000000000000000", 10018 => "0000000000000000", 10019 => "0000000000000000", 10020 => "0000000000000000", 10021 => "0000000000000000", 10022 => "0000000000000000", 10023 => "0000000000000000", 10024 => "0000000000000000", 10025 => "0000000000000000", 10026 => "0000000000000000", 10027 => "0000000000000000", 10028 => "0000000000000000", 10029 => "0000000000000000", 10030 => "0000000000000000", 10031 => "0000000000000000", 10032 => "0000000000000000", 10033 => "0000000000000000", 10034 => "0000000000000000", 10035 => "0000000000000000", 10036 => "0000000000000000", 10037 => "0000000000000000", 10038 => "0000000000000000", 10039 => "0000000000000000", 10040 => "0000000000000000", 10041 => "0000000000000000", 10042 => "0000000000000000", 10043 => "0000000000000000", 10044 => "0000000000000000", 10045 => "0000000000000000", 10046 => "0000000000000000", 10047 => "0000000000000000", 10048 => "0000000000000000", 10049 => "0000000000000000", 10050 => "0000000000000000", 10051 => "0000000000000000", 10052 => "0000000000000000", 10053 => "0000000000000000", 10054 => "0000000000000000", 10055 => "0000000000000000", 10056 => "0000000000000000", 10057 => "0000000000000000", 10058 => "0000000000000000", 10059 => "0000000000000000", 10060 => "0000000000000000", 10061 => "0000000000000000", 10062 => "0000000000000000", 10063 => "0000000000000000", 10064 => "0000000000000000", 10065 => "0000000000000000", 10066 => "0000000000000000", 10067 => "0000000000000000", 10068 => "0000000000000000", 10069 => "0000000000000000", 10070 => "0000000000000000", 10071 => "0000000000000000", 10072 => "0000000000000000", 10073 => "0000000000000000", 10074 => "0000000000000000", 10075 => "0000000000000000", 10076 => "0000000000000000", 10077 => "0000000000000000", 10078 => "0000000000000000", 10079 => "0000000000000000", 10080 => "0000000000000000", 10081 => "0000000000000000", 10082 => "0000000000000000", 10083 => "0000000000000000", 10084 => "0000000000000000", 10085 => "0000000000000000", 10086 => "0000000000000000", 10087 => "0000000000000000", 10088 => "0000000000000000", 10089 => "0000000000000000", 10090 => "0000000000000000", 10091 => "0000000000000000", 10092 => "0000000000000000", 10093 => "0000000000000000", 10094 => "0000000000000000", 10095 => "0000000000000000", 10096 => "0000000000000000", 10097 => "0000000000000000", 10098 => "0000000000000000", 10099 => "0000000000000000", 10100 => "0000000000000000", 10101 => "0000000000000000", 10102 => "0000000000000000", 10103 => "0000000000000000", 10104 => "0000000000000000", 10105 => "0000000000000000", 10106 => "0000000000000000", 10107 => "0000000000000000", 10108 => "0000000000000000", 10109 => "0000000000000000", 10110 => "0000000000000000", 10111 => "0000000000000000", 10112 => "0000000000000000", 10113 => "0000000000000000", 10114 => "0000000000000000", 10115 => "0000000000000000", 10116 => "0000000000000000", 10117 => "0000000000000000", 10118 => "0000000000000000", 10119 => "0000000000000000", 10120 => "0000000000000000", 10121 => "0000000000000000", 10122 => "0000000000000000", 10123 => "0000000000000000", 10124 => "0000000000000000", 10125 => "0000000000000000", 10126 => "0000000000000000", 10127 => "0000000000000000", 10128 => "0000000000000000", 10129 => "0000000000000000", 10130 => "0000000000000000", 10131 => "0000000000000000", 10132 => "0000000000000000", 10133 => "0000000000000000", 10134 => "0000000000000000", 10135 => "0000000000000000", 10136 => "0000000000000000", 10137 => "0000000000000000", 10138 => "0000000000000000", 10139 => "0000000000000000", 10140 => "0000000000000000", 10141 => "0000000000000000", 10142 => "0000000000000000", 10143 => "0000000000000000", 10144 => "0000000000000000", 10145 => "0000000000000000", 10146 => "0000000000000000", 10147 => "0000000000000000", 10148 => "0000000000000000", 10149 => "0000000000000000", 10150 => "0000000000000000", 10151 => "0000000000000000", 10152 => "0000000000000000", 10153 => "0000000000000000", 10154 => "0000000000000000", 10155 => "0000000000000000", 10156 => "0000000000000000", 10157 => "0000000000000000", 10158 => "0000000000000000", 10159 => "0000000000000000", 10160 => "0000000000000000", 10161 => "0000000000000000", 10162 => "0000000000000000", 10163 => "0000000000000000", 10164 => "0000000000000000", 10165 => "0000000000000000", 10166 => "0000000000000000", 10167 => "0000000000000000", 10168 => "0000000000000000", 10169 => "0000000000000000", 10170 => "0000000000000000", 10171 => "0000000000000000", 10172 => "0000000000000000", 10173 => "0000000000000000", 10174 => "0000000000000000", 10175 => "0000000000000000", 10176 => "0000000000000000", 10177 => "0000000000000000", 10178 => "0000000000000000", 10179 => "0000000000000000", 10180 => "0000000000000000", 10181 => "0000000000000000", 10182 => "0000000000000000", 10183 => "0000000000000000", 10184 => "0000000000000000", 10185 => "0000000000000000", 10186 => "0000000000000000", 10187 => "0000000000000000", 10188 => "0000000000000000", 10189 => "0000000000000000", 10190 => "0000000000000000", 10191 => "0000000000000000", 10192 => "0000000000000000", 10193 => "0000000000000000", 10194 => "0000000000000000", 10195 => "0000000000000000", 10196 => "0000000000000000", 10197 => "0000000000000000", 10198 => "0000000000000000", 10199 => "0000000000000000", 10200 => "0000000000000000", 10201 => "0000000000000000", 10202 => "0000000000000000", 10203 => "0000000000000000", 10204 => "0000000000000000", 10205 => "0000000000000000", 10206 => "0000000000000000", 10207 => "0000000000000000", 10208 => "0000000000000000", 10209 => "0000000000000000", 10210 => "0000000000000000", 10211 => "0000000000000000", 10212 => "0000000000000000", 10213 => "0000000000000000", 10214 => "0000000000000000", 10215 => "0000000000000000", 10216 => "0000000000000000", 10217 => "0000000000000000", 10218 => "0000000000000000", 10219 => "0000000000000000", 10220 => "0000000000000000", 10221 => "0000000000000000", 10222 => "0000000000000000", 10223 => "0000000000000000", 10224 => "0000000000000000", 10225 => "0000000000000000", 10226 => "0000000000000000", 10227 => "0000000000000000", 10228 => "0000000000000000", 10229 => "0000000000000000", 10230 => "0000000000000000", 10231 => "0000000000000000", 10232 => "0000000000000000", 10233 => "0000000000000000", 10234 => "0000000000000000", 10235 => "0000000000000000", 10236 => "0000000000000000", 10237 => "0000000000000000", 10238 => "0000000000000000", 10239 => "0000000000000000", 10240 => "0000000000000000", 10241 => "0000000000000000", 10242 => "0000000000000000", 10243 => "0000000000000000", 10244 => "0000000000000000", 10245 => "0000000000000000", 10246 => "0000000000000000", 10247 => "0000000000000000", 10248 => "0000000000000000", 10249 => "0000000000000000", 10250 => "0000000000000000", 10251 => "0000000000000000", 10252 => "0000000000000000", 10253 => "0000000000000000", 10254 => "0000000000000000", 10255 => "0000000000000000", 10256 => "0000000000000000", 10257 => "0000000000000000", 10258 => "0000000000000000", 10259 => "0000000000000000", 10260 => "0000000000000000", 10261 => "0000000000000000", 10262 => "0000000000000000", 10263 => "0000000000000000", 10264 => "0000000000000000", 10265 => "0000000000000000", 10266 => "0000000000000000", 10267 => "0000000000000000", 10268 => "0000000000000000", 10269 => "0000000000000000", 10270 => "0000000000000000", 10271 => "0000000000000000", 10272 => "0000000000000000", 10273 => "0000000000000000", 10274 => "0000000000000000", 10275 => "0000000000000000", 10276 => "0000000000000000", 10277 => "0000000000000000", 10278 => "0000000000000000", 10279 => "0000000000000000", 10280 => "0000000000000000", 10281 => "0000000000000000", 10282 => "0000000000000000", 10283 => "0000000000000000", 10284 => "0000000000000000", 10285 => "0000000000000000", 10286 => "0000000000000000", 10287 => "0000000000000000", 10288 => "0000000000000000", 10289 => "0000000000000000", 10290 => "0000000000000000", 10291 => "0000000000000000", 10292 => "0000000000000000", 10293 => "0000000000000000", 10294 => "0000000000000000", 10295 => "0000000000000000", 10296 => "0000000000000000", 10297 => "0000000000000000", 10298 => "0000000000000000", 10299 => "0000000000000000", 10300 => "0000000000000000", 10301 => "0000000000000000", 10302 => "0000000000000000", 10303 => "0000000000000000", 10304 => "0000000000000000", 10305 => "0000000000000000", 10306 => "0000000000000000", 10307 => "0000000000000000", 10308 => "0000000000000000", 10309 => "0000000000000000", 10310 => "0000000000000000", 10311 => "0000000000000000", 10312 => "0000000000000000", 10313 => "0000000000000000", 10314 => "0000000000000000", 10315 => "0000000000000000", 10316 => "0000000000000000", 10317 => "0000000000000000", 10318 => "0000000000000000", 10319 => "0000000000000000", 10320 => "0000000000000000", 10321 => "0000000000000000", 10322 => "0000000000000000", 10323 => "0000000000000000", 10324 => "0000000000000000", 10325 => "0000000000000000", 10326 => "0000000000000000", 10327 => "0000000000000000", 10328 => "0000000000000000", 10329 => "0000000000000000", 10330 => "0000000000000000", 10331 => "0000000000000000", 10332 => "0000000000000000", 10333 => "0000000000000000", 10334 => "0000000000000000", 10335 => "0000000000000000", 10336 => "0000000000000000", 10337 => "0000000000000000", 10338 => "0000000000000000", 10339 => "0000000000000000", 10340 => "0000000000000000", 10341 => "0000000000000000", 10342 => "0000000000000000", 10343 => "0000000000000000", 10344 => "0000000000000000", 10345 => "0000000000000000", 10346 => "0000000000000000", 10347 => "0000000000000000", 10348 => "0000000000000000", 10349 => "0000000000000000", 10350 => "0000000000000000", 10351 => "0000000000000000", 10352 => "0000000000000000", 10353 => "0000000000000000", 10354 => "0000000000000000", 10355 => "0000000000000000", 10356 => "0000000000000000", 10357 => "0000000000000000", 10358 => "0000000000000000", 10359 => "0000000000000000", 10360 => "0000000000000000", 10361 => "0000000000000000", 10362 => "0000000000000000", 10363 => "0000000000000000", 10364 => "0000000000000000", 10365 => "0000000000000000", 10366 => "0000000000000000", 10367 => "0000000000000000", 10368 => "0000000000000000", 10369 => "0000000000000000", 10370 => "0000000000000000", 10371 => "0000000000000000", 10372 => "0000000000000000", 10373 => "0000000000000000", 10374 => "0000000000000000", 10375 => "0000000000000000", 10376 => "0000000000000000", 10377 => "0000000000000000", 10378 => "0000000000000000", 10379 => "0000000000000000", 10380 => "0000000000000000", 10381 => "0000000000000000", 10382 => "0000000000000000", 10383 => "0000000000000000", 10384 => "0000000000000000", 10385 => "0000000000000000", 10386 => "0000000000000000", 10387 => "0000000000000000", 10388 => "0000000000000000", 10389 => "0000000000000000", 10390 => "0000000000000000", 10391 => "0000000000000000", 10392 => "0000000000000000", 10393 => "0000000000000000", 10394 => "0000000000000000", 10395 => "0000000000000000", 10396 => "0000000000000000", 10397 => "0000000000000000", 10398 => "0000000000000000", 10399 => "0000000000000000", 10400 => "0000000000000000", 10401 => "0000000000000000", 10402 => "0000000000000000", 10403 => "0000000000000000", 10404 => "0000000000000000", 10405 => "0000000000000000", 10406 => "0000000000000000", 10407 => "0000000000000000", 10408 => "0000000000000000", 10409 => "0000000000000000", 10410 => "0000000000000000", 10411 => "0000000000000000", 10412 => "0000000000000000", 10413 => "0000000000000000", 10414 => "0000000000000000", 10415 => "0000000000000000", 10416 => "0000000000000000", 10417 => "0000000000000000", 10418 => "0000000000000000", 10419 => "0000000000000000", 10420 => "0000000000000000", 10421 => "0000000000000000", 10422 => "0000000000000000", 10423 => "0000000000000000", 10424 => "0000000000000000", 10425 => "0000000000000000", 10426 => "0000000000000000", 10427 => "0000000000000000", 10428 => "0000000000000000", 10429 => "0000000000000000", 10430 => "0000000000000000", 10431 => "0000000000000000", 10432 => "0000000000000000", 10433 => "0000000000000000", 10434 => "0000000000000000", 10435 => "0000000000000000", 10436 => "0000000000000000", 10437 => "0000000000000000", 10438 => "0000000000000000", 10439 => "0000000000000000", 10440 => "0000000000000000", 10441 => "0000000000000000", 10442 => "0000000000000000", 10443 => "0000000000000000", 10444 => "0000000000000000", 10445 => "0000000000000000", 10446 => "0000000000000000", 10447 => "0000000000000000", 10448 => "0000000000000000", 10449 => "0000000000000000", 10450 => "0000000000000000", 10451 => "0000000000000000", 10452 => "0000000000000000", 10453 => "0000000000000000", 10454 => "0000000000000000", 10455 => "0000000000000000", 10456 => "0000000000000000", 10457 => "0000000000000000", 10458 => "0000000000000000", 10459 => "0000000000000000", 10460 => "0000000000000000", 10461 => "0000000000000000", 10462 => "0000000000000000", 10463 => "0000000000000000", 10464 => "0000000000000000", 10465 => "0000000000000000", 10466 => "0000000000000000", 10467 => "0000000000000000", 10468 => "0000000000000000", 10469 => "0000000000000000", 10470 => "0000000000000000", 10471 => "0000000000000000", 10472 => "0000000000000000", 10473 => "0000000000000000", 10474 => "0000000000000000", 10475 => "0000000000000000", 10476 => "0000000000000000", 10477 => "0000000000000000", 10478 => "0000000000000000", 10479 => "0000000000000000", 10480 => "0000000000000000", 10481 => "0000000000000000", 10482 => "0000000000000000", 10483 => "0000000000000000", 10484 => "0000000000000000", 10485 => "0000000000000000", 10486 => "0000000000000000", 10487 => "0000000000000000", 10488 => "0000000000000000", 10489 => "0000000000000000", 10490 => "0000000000000000", 10491 => "0000000000000000", 10492 => "0000000000000000", 10493 => "0000000000000000", 10494 => "0000000000000000", 10495 => "0000000000000000", 10496 => "0000000000000000", 10497 => "0000000000000000", 10498 => "0000000000000000", 10499 => "0000000000000000", 10500 => "0000000000000000", 10501 => "0000000000000000", 10502 => "0000000000000000", 10503 => "0000000000000000", 10504 => "0000000000000000", 10505 => "0000000000000000", 10506 => "0000000000000000", 10507 => "0000000000000000", 10508 => "0000000000000000", 10509 => "0000000000000000", 10510 => "0000000000000000", 10511 => "0000000000000000", 10512 => "0000000000000000", 10513 => "0000000000000000", 10514 => "0000000000000000", 10515 => "0000000000000000", 10516 => "0000000000000000", 10517 => "0000000000000000", 10518 => "0000000000000000", 10519 => "0000000000000000", 10520 => "0000000000000000", 10521 => "0000000000000000", 10522 => "0000000000000000", 10523 => "0000000000000000", 10524 => "0000000000000000", 10525 => "0000000000000000", 10526 => "0000000000000000", 10527 => "0000000000000000", 10528 => "0000000000000000", 10529 => "0000000000000000", 10530 => "0000000000000000", 10531 => "0000000000000000", 10532 => "0000000000000000", 10533 => "0000000000000000", 10534 => "0000000000000000", 10535 => "0000000000000000", 10536 => "0000000000000000", 10537 => "0000000000000000", 10538 => "0000000000000000", 10539 => "0000000000000000", 10540 => "0000000000000000", 10541 => "0000000000000000", 10542 => "0000000000000000", 10543 => "0000000000000000", 10544 => "0000000000000000", 10545 => "0000000000000000", 10546 => "0000000000000000", 10547 => "0000000000000000", 10548 => "0000000000000000", 10549 => "0000000000000000", 10550 => "0000000000000000", 10551 => "0000000000000000", 10552 => "0000000000000000", 10553 => "0000000000000000", 10554 => "0000000000000000", 10555 => "0000000000000000", 10556 => "0000000000000000", 10557 => "0000000000000000", 10558 => "0000000000000000", 10559 => "0000000000000000", 10560 => "0000000000000000", 10561 => "0000000000000000", 10562 => "0000000000000000", 10563 => "0000000000000000", 10564 => "0000000000000000", 10565 => "0000000000000000", 10566 => "0000000000000000", 10567 => "0000000000000000", 10568 => "0000000000000000", 10569 => "0000000000000000", 10570 => "0000000000000000", 10571 => "0000000000000000", 10572 => "0000000000000000", 10573 => "0000000000000000", 10574 => "0000000000000000", 10575 => "0000000000000000", 10576 => "0000000000000000", 10577 => "0000000000000000", 10578 => "0000000000000000", 10579 => "0000000000000000", 10580 => "0000000000000000", 10581 => "0000000000000000", 10582 => "0000000000000000", 10583 => "0000000000000000", 10584 => "0000000000000000", 10585 => "0000000000000000", 10586 => "0000000000000000", 10587 => "0000000000000000", 10588 => "0000000000000000", 10589 => "0000000000000000", 10590 => "0000000000000000", 10591 => "0000000000000000", 10592 => "0000000000000000", 10593 => "0000000000000000", 10594 => "0000000000000000", 10595 => "0000000000000000", 10596 => "0000000000000000", 10597 => "0000000000000000", 10598 => "0000000000000000", 10599 => "0000000000000000", 10600 => "0000000000000000", 10601 => "0000000000000000", 10602 => "0000000000000000", 10603 => "0000000000000000", 10604 => "0000000000000000", 10605 => "0000000000000000", 10606 => "0000000000000000", 10607 => "0000000000000000", 10608 => "0000000000000000", 10609 => "0000000000000000", 10610 => "0000000000000000", 10611 => "0000000000000000", 10612 => "0000000000000000", 10613 => "0000000000000000", 10614 => "0000000000000000", 10615 => "0000000000000000", 10616 => "0000000000000000", 10617 => "0000000000000000", 10618 => "0000000000000000", 10619 => "0000000000000000", 10620 => "0000000000000000", 10621 => "0000000000000000", 10622 => "0000000000000000", 10623 => "0000000000000000", 10624 => "0000000000000000", 10625 => "0000000000000000", 10626 => "0000000000000000", 10627 => "0000000000000000", 10628 => "0000000000000000", 10629 => "0000000000000000", 10630 => "0000000000000000", 10631 => "0000000000000000", 10632 => "0000000000000000", 10633 => "0000000000000000", 10634 => "0000000000000000", 10635 => "0000000000000000", 10636 => "0000000000000000", 10637 => "0000000000000000", 10638 => "0000000000000000", 10639 => "0000000000000000", 10640 => "0000000000000000", 10641 => "0000000000000000", 10642 => "0000000000000000", 10643 => "0000000000000000", 10644 => "0000000000000000", 10645 => "0000000000000000", 10646 => "0000000000000000", 10647 => "0000000000000000", 10648 => "0000000000000000", 10649 => "0000000000000000", 10650 => "0000000000000000", 10651 => "0000000000000000", 10652 => "0000000000000000", 10653 => "0000000000000000", 10654 => "0000000000000000", 10655 => "0000000000000000", 10656 => "0000000000000000", 10657 => "0000000000000000", 10658 => "0000000000000000", 10659 => "0000000000000000", 10660 => "0000000000000000", 10661 => "0000000000000000", 10662 => "0000000000000000", 10663 => "0000000000000000", 10664 => "0000000000000000", 10665 => "0000000000000000", 10666 => "0000000000000000", 10667 => "0000000000000000", 10668 => "0000000000000000", 10669 => "0000000000000000", 10670 => "0000000000000000", 10671 => "0000000000000000", 10672 => "0000000000000000", 10673 => "0000000000000000", 10674 => "0000000000000000", 10675 => "0000000000000000", 10676 => "0000000000000000", 10677 => "0000000000000000", 10678 => "0000000000000000", 10679 => "0000000000000000", 10680 => "0000000000000000", 10681 => "0000000000000000", 10682 => "0000000000000000", 10683 => "0000000000000000", 10684 => "0000000000000000", 10685 => "0000000000000000", 10686 => "0000000000000000", 10687 => "0000000000000000", 10688 => "0000000000000000", 10689 => "0000000000000000", 10690 => "0000000000000000", 10691 => "0000000000000000", 10692 => "0000000000000000", 10693 => "0000000000000000", 10694 => "0000000000000000", 10695 => "0000000000000000", 10696 => "0000000000000000", 10697 => "0000000000000000", 10698 => "0000000000000000", 10699 => "0000000000000000", 10700 => "0000000000000000", 10701 => "0000000000000000", 10702 => "0000000000000000", 10703 => "0000000000000000", 10704 => "0000000000000000", 10705 => "0000000000000000", 10706 => "0000000000000000", 10707 => "0000000000000000", 10708 => "0000000000000000", 10709 => "0000000000000000", 10710 => "0000000000000000", 10711 => "0000000000000000", 10712 => "0000000000000000", 10713 => "0000000000000000", 10714 => "0000000000000000", 10715 => "0000000000000000", 10716 => "0000000000000000", 10717 => "0000000000000000", 10718 => "0000000000000000", 10719 => "0000000000000000", 10720 => "0000000000000000", 10721 => "0000000000000000", 10722 => "0000000000000000", 10723 => "0000000000000000", 10724 => "0000000000000000", 10725 => "0000000000000000", 10726 => "0000000000000000", 10727 => "0000000000000000", 10728 => "0000000000000000", 10729 => "0000000000000000", 10730 => "0000000000000000", 10731 => "0000000000000000", 10732 => "0000000000000000", 10733 => "0000000000000000", 10734 => "0000000000000000", 10735 => "0000000000000000", 10736 => "0000000000000000", 10737 => "0000000000000000", 10738 => "0000000000000000", 10739 => "0000000000000000", 10740 => "0000000000000000", 10741 => "0000000000000000", 10742 => "0000000000000000", 10743 => "0000000000000000", 10744 => "0000000000000000", 10745 => "0000000000000000", 10746 => "0000000000000000", 10747 => "0000000000000000", 10748 => "0000000000000000", 10749 => "0000000000000000", 10750 => "0000000000000000", 10751 => "0000000000000000", 10752 => "0000000000000000", 10753 => "0000000000000000", 10754 => "0000000000000000", 10755 => "0000000000000000", 10756 => "0000000000000000", 10757 => "0000000000000000", 10758 => "0000000000000000", 10759 => "0000000000000000", 10760 => "0000000000000000", 10761 => "0000000000000000", 10762 => "0000000000000000", 10763 => "0000000000000000", 10764 => "0000000000000000", 10765 => "0000000000000000", 10766 => "0000000000000000", 10767 => "0000000000000000", 10768 => "0000000000000000", 10769 => "0000000000000000", 10770 => "0000000000000000", 10771 => "0000000000000000", 10772 => "0000000000000000", 10773 => "0000000000000000", 10774 => "0000000000000000", 10775 => "0000000000000000", 10776 => "0000000000000000", 10777 => "0000000000000000", 10778 => "0000000000000000", 10779 => "0000000000000000", 10780 => "0000000000000000", 10781 => "0000000000000000", 10782 => "0000000000000000", 10783 => "0000000000000000", 10784 => "0000000000000000", 10785 => "0000000000000000", 10786 => "0000000000000000", 10787 => "0000000000000000", 10788 => "0000000000000000", 10789 => "0000000000000000", 10790 => "0000000000000000", 10791 => "0000000000000000", 10792 => "0000000000000000", 10793 => "0000000000000000", 10794 => "0000000000000000", 10795 => "0000000000000000", 10796 => "0000000000000000", 10797 => "0000000000000000", 10798 => "0000000000000000", 10799 => "0000000000000000", 10800 => "0000000000000000", 10801 => "0000000000000000", 10802 => "0000000000000000", 10803 => "0000000000000000", 10804 => "0000000000000000", 10805 => "0000000000000000", 10806 => "0000000000000000", 10807 => "0000000000000000", 10808 => "0000000000000000", 10809 => "0000000000000000", 10810 => "0000000000000000", 10811 => "0000000000000000", 10812 => "0000000000000000", 10813 => "0000000000000000", 10814 => "0000000000000000", 10815 => "0000000000000000", 10816 => "0000000000000000", 10817 => "0000000000000000", 10818 => "0000000000000000", 10819 => "0000000000000000", 10820 => "0000000000000000", 10821 => "0000000000000000", 10822 => "0000000000000000", 10823 => "0000000000000000", 10824 => "0000000000000000", 10825 => "0000000000000000", 10826 => "0000000000000000", 10827 => "0000000000000000", 10828 => "0000000000000000", 10829 => "0000000000000000", 10830 => "0000000000000000", 10831 => "0000000000000000", 10832 => "0000000000000000", 10833 => "0000000000000000", 10834 => "0000000000000000", 10835 => "0000000000000000", 10836 => "0000000000000000", 10837 => "0000000000000000", 10838 => "0000000000000000", 10839 => "0000000000000000", 10840 => "0000000000000000", 10841 => "0000000000000000", 10842 => "0000000000000000", 10843 => "0000000000000000", 10844 => "0000000000000000", 10845 => "0000000000000000", 10846 => "0000000000000000", 10847 => "0000000000000000", 10848 => "0000000000000000", 10849 => "0000000000000000", 10850 => "0000000000000000", 10851 => "0000000000000000", 10852 => "0000000000000000", 10853 => "0000000000000000", 10854 => "0000000000000000", 10855 => "0000000000000000", 10856 => "0000000000000000", 10857 => "0000000000000000", 10858 => "0000000000000000", 10859 => "0000000000000000", 10860 => "0000000000000000", 10861 => "0000000000000000", 10862 => "0000000000000000", 10863 => "0000000000000000", 10864 => "0000000000000000", 10865 => "0000000000000000", 10866 => "0000000000000000", 10867 => "0000000000000000", 10868 => "0000000000000000", 10869 => "0000000000000000", 10870 => "0000000000000000", 10871 => "0000000000000000", 10872 => "0000000000000000", 10873 => "0000000000000000", 10874 => "0000000000000000", 10875 => "0000000000000000", 10876 => "0000000000000000", 10877 => "0000000000000000", 10878 => "0000000000000000", 10879 => "0000000000000000", 10880 => "0000000000000000", 10881 => "0000000000000000", 10882 => "0000000000000000", 10883 => "0000000000000000", 10884 => "0000000000000000", 10885 => "0000000000000000", 10886 => "0000000000000000", 10887 => "0000000000000000", 10888 => "0000000000000000", 10889 => "0000000000000000", 10890 => "0000000000000000", 10891 => "0000000000000000", 10892 => "0000000000000000", 10893 => "0000000000000000", 10894 => "0000000000000000", 10895 => "0000000000000000", 10896 => "0000000000000000", 10897 => "0000000000000000", 10898 => "0000000000000000", 10899 => "0000000000000000", 10900 => "0000000000000000", 10901 => "0000000000000000", 10902 => "0000000000000000", 10903 => "0000000000000000", 10904 => "0000000000000000", 10905 => "0000000000000000", 10906 => "0000000000000000", 10907 => "0000000000000000", 10908 => "0000000000000000", 10909 => "0000000000000000", 10910 => "0000000000000000", 10911 => "0000000000000000", 10912 => "0000000000000000", 10913 => "0000000000000000", 10914 => "0000000000000000", 10915 => "0000000000000000", 10916 => "0000000000000000", 10917 => "0000000000000000", 10918 => "0000000000000000", 10919 => "0000000000000000", 10920 => "0000000000000000", 10921 => "0000000000000000", 10922 => "0000000000000000", 10923 => "0000000000000000", 10924 => "0000000000000000", 10925 => "0000000000000000", 10926 => "0000000000000000", 10927 => "0000000000000000", 10928 => "0000000000000000", 10929 => "0000000000000000", 10930 => "0000000000000000", 10931 => "0000000000000000", 10932 => "0000000000000000", 10933 => "0000000000000000", 10934 => "0000000000000000", 10935 => "0000000000000000", 10936 => "0000000000000000", 10937 => "0000000000000000", 10938 => "0000000000000000", 10939 => "0000000000000000", 10940 => "0000000000000000", 10941 => "0000000000000000", 10942 => "0000000000000000", 10943 => "0000000000000000", 10944 => "0000000000000000", 10945 => "0000000000000000", 10946 => "0000000000000000", 10947 => "0000000000000000", 10948 => "0000000000000000", 10949 => "0000000000000000", 10950 => "0000000000000000", 10951 => "0000000000000000", 10952 => "0000000000000000", 10953 => "0000000000000000", 10954 => "0000000000000000", 10955 => "0000000000000000", 10956 => "0000000000000000", 10957 => "0000000000000000", 10958 => "0000000000000000", 10959 => "0000000000000000", 10960 => "0000000000000000", 10961 => "0000000000000000", 10962 => "0000000000000000", 10963 => "0000000000000000", 10964 => "0000000000000000", 10965 => "0000000000000000", 10966 => "0000000000000000", 10967 => "0000000000000000", 10968 => "0000000000000000", 10969 => "0000000000000000", 10970 => "0000000000000000", 10971 => "0000000000000000", 10972 => "0000000000000000", 10973 => "0000000000000000", 10974 => "0000000000000000", 10975 => "0000000000000000", 10976 => "0000000000000000", 10977 => "0000000000000000", 10978 => "0000000000000000", 10979 => "0000000000000000", 10980 => "0000000000000000", 10981 => "0000000000000000", 10982 => "0000000000000000", 10983 => "0000000000000000", 10984 => "0000000000000000", 10985 => "0000000000000000", 10986 => "0000000000000000", 10987 => "0000000000000000", 10988 => "0000000000000000", 10989 => "0000000000000000", 10990 => "0000000000000000", 10991 => "0000000000000000", 10992 => "0000000000000000", 10993 => "0000000000000000", 10994 => "0000000000000000", 10995 => "0000000000000000", 10996 => "0000000000000000", 10997 => "0000000000000000", 10998 => "0000000000000000", 10999 => "0000000000000000", 11000 => "0000000000000000", 11001 => "0000000000000000", 11002 => "0000000000000000", 11003 => "0000000000000000", 11004 => "0000000000000000", 11005 => "0000000000000000", 11006 => "0000000000000000", 11007 => "0000000000000000", 11008 => "0000000000000000", 11009 => "0000000000000000", 11010 => "0000000000000000", 11011 => "0000000000000000", 11012 => "0000000000000000", 11013 => "0000000000000000", 11014 => "0000000000000000", 11015 => "0000000000000000", 11016 => "0000000000000000", 11017 => "0000000000000000", 11018 => "0000000000000000", 11019 => "0000000000000000", 11020 => "0000000000000000", 11021 => "0000000000000000", 11022 => "0000000000000000", 11023 => "0000000000000000", 11024 => "0000000000000000", 11025 => "0000000000000000", 11026 => "0000000000000000", 11027 => "0000000000000000", 11028 => "0000000000000000", 11029 => "0000000000000000", 11030 => "0000000000000000", 11031 => "0000000000000000", 11032 => "0000000000000000", 11033 => "0000000000000000", 11034 => "0000000000000000", 11035 => "0000000000000000", 11036 => "0000000000000000", 11037 => "0000000000000000", 11038 => "0000000000000000", 11039 => "0000000000000000", 11040 => "0000000000000000", 11041 => "0000000000000000", 11042 => "0000000000000000", 11043 => "0000000000000000", 11044 => "0000000000000000", 11045 => "0000000000000000", 11046 => "0000000000000000", 11047 => "0000000000000000", 11048 => "0000000000000000", 11049 => "0000000000000000", 11050 => "0000000000000000", 11051 => "0000000000000000", 11052 => "0000000000000000", 11053 => "0000000000000000", 11054 => "0000000000000000", 11055 => "0000000000000000", 11056 => "0000000000000000", 11057 => "0000000000000000", 11058 => "0000000000000000", 11059 => "0000000000000000", 11060 => "0000000000000000", 11061 => "0000000000000000", 11062 => "0000000000000000", 11063 => "0000000000000000", 11064 => "0000000000000000", 11065 => "0000000000000000", 11066 => "0000000000000000", 11067 => "0000000000000000", 11068 => "0000000000000000", 11069 => "0000000000000000", 11070 => "0000000000000000", 11071 => "0000000000000000", 11072 => "0000000000000000", 11073 => "0000000000000000", 11074 => "0000000000000000", 11075 => "0000000000000000", 11076 => "0000000000000000", 11077 => "0000000000000000", 11078 => "0000000000000000", 11079 => "0000000000000000", 11080 => "0000000000000000", 11081 => "0000000000000000", 11082 => "0000000000000000", 11083 => "0000000000000000", 11084 => "0000000000000000", 11085 => "0000000000000000", 11086 => "0000000000000000", 11087 => "0000000000000000", 11088 => "0000000000000000", 11089 => "0000000000000000", 11090 => "0000000000000000", 11091 => "0000000000000000", 11092 => "0000000000000000", 11093 => "0000000000000000", 11094 => "0000000000000000", 11095 => "0000000000000000", 11096 => "0000000000000000", 11097 => "0000000000000000", 11098 => "0000000000000000", 11099 => "0000000000000000", 11100 => "0000000000000000", 11101 => "0000000000000000", 11102 => "0000000000000000", 11103 => "0000000000000000", 11104 => "0000000000000000", 11105 => "0000000000000000", 11106 => "0000000000000000", 11107 => "0000000000000000", 11108 => "0000000000000000", 11109 => "0000000000000000", 11110 => "0000000000000000", 11111 => "0000000000000000", 11112 => "0000000000000000", 11113 => "0000000000000000", 11114 => "0000000000000000", 11115 => "0000000000000000", 11116 => "0000000000000000", 11117 => "0000000000000000", 11118 => "0000000000000000", 11119 => "0000000000000000", 11120 => "0000000000000000", 11121 => "0000000000000000", 11122 => "0000000000000000", 11123 => "0000000000000000", 11124 => "0000000000000000", 11125 => "0000000000000000", 11126 => "0000000000000000", 11127 => "0000000000000000", 11128 => "0000000000000000", 11129 => "0000000000000000", 11130 => "0000000000000000", 11131 => "0000000000000000", 11132 => "0000000000000000", 11133 => "0000000000000000", 11134 => "0000000000000000", 11135 => "0000000000000000", 11136 => "0000000000000000", 11137 => "0000000000000000", 11138 => "0000000000000000", 11139 => "0000000000000000", 11140 => "0000000000000000", 11141 => "0000000000000000", 11142 => "0000000000000000", 11143 => "0000000000000000", 11144 => "0000000000000000", 11145 => "0000000000000000", 11146 => "0000000000000000", 11147 => "0000000000000000", 11148 => "0000000000000000", 11149 => "0000000000000000", 11150 => "0000000000000000", 11151 => "0000000000000000", 11152 => "0000000000000000", 11153 => "0000000000000000", 11154 => "0000000000000000", 11155 => "0000000000000000", 11156 => "0000000000000000", 11157 => "0000000000000000", 11158 => "0000000000000000", 11159 => "0000000000000000", 11160 => "0000000000000000", 11161 => "0000000000000000", 11162 => "0000000000000000", 11163 => "0000000000000000", 11164 => "0000000000000000", 11165 => "0000000000000000", 11166 => "0000000000000000", 11167 => "0000000000000000", 11168 => "0000000000000000", 11169 => "0000000000000000", 11170 => "0000000000000000", 11171 => "0000000000000000", 11172 => "0000000000000000", 11173 => "0000000000000000", 11174 => "0000000000000000", 11175 => "0000000000000000", 11176 => "0000000000000000", 11177 => "0000000000000000", 11178 => "0000000000000000", 11179 => "0000000000000000", 11180 => "0000000000000000", 11181 => "0000000000000000", 11182 => "0000000000000000", 11183 => "0000000000000000", 11184 => "0000000000000000", 11185 => "0000000000000000", 11186 => "0000000000000000", 11187 => "0000000000000000", 11188 => "0000000000000000", 11189 => "0000000000000000", 11190 => "0000000000000000", 11191 => "0000000000000000", 11192 => "0000000000000000", 11193 => "0000000000000000", 11194 => "0000000000000000", 11195 => "0000000000000000", 11196 => "0000000000000000", 11197 => "0000000000000000", 11198 => "0000000000000000", 11199 => "0000000000000000", 11200 => "0000000000000000", 11201 => "0000000000000000", 11202 => "0000000000000000", 11203 => "0000000000000000", 11204 => "0000000000000000", 11205 => "0000000000000000", 11206 => "0000000000000000", 11207 => "0000000000000000", 11208 => "0000000000000000", 11209 => "0000000000000000", 11210 => "0000000000000000", 11211 => "0000000000000000", 11212 => "0000000000000000", 11213 => "0000000000000000", 11214 => "0000000000000000", 11215 => "0000000000000000", 11216 => "0000000000000000", 11217 => "0000000000000000", 11218 => "0000000000000000", 11219 => "0000000000000000", 11220 => "0000000000000000", 11221 => "0000000000000000", 11222 => "0000000000000000", 11223 => "0000000000000000", 11224 => "0000000000000000", 11225 => "0000000000000000", 11226 => "0000000000000000", 11227 => "0000000000000000", 11228 => "0000000000000000", 11229 => "0000000000000000", 11230 => "0000000000000000", 11231 => "0000000000000000", 11232 => "0000000000000000", 11233 => "0000000000000000", 11234 => "0000000000000000", 11235 => "0000000000000000", 11236 => "0000000000000000", 11237 => "0000000000000000", 11238 => "0000000000000000", 11239 => "0000000000000000", 11240 => "0000000000000000", 11241 => "0000000000000000", 11242 => "0000000000000000", 11243 => "0000000000000000", 11244 => "0000000000000000", 11245 => "0000000000000000", 11246 => "0000000000000000", 11247 => "0000000000000000", 11248 => "0000000000000000", 11249 => "0000000000000000", 11250 => "0000000000000000", 11251 => "0000000000000000", 11252 => "0000000000000000", 11253 => "0000000000000000", 11254 => "0000000000000000", 11255 => "0000000000000000", 11256 => "0000000000000000", 11257 => "0000000000000000", 11258 => "0000000000000000", 11259 => "0000000000000000", 11260 => "0000000000000000", 11261 => "0000000000000000", 11262 => "0000000000000000", 11263 => "0000000000000000", 11264 => "0000000000000000", 11265 => "0000000000000000", 11266 => "0000000000000000", 11267 => "0000000000000000", 11268 => "0000000000000000", 11269 => "0000000000000000", 11270 => "0000000000000000", 11271 => "0000000000000000", 11272 => "0000000000000000", 11273 => "0000000000000000", 11274 => "0000000000000000", 11275 => "0000000000000000", 11276 => "0000000000000000", 11277 => "0000000000000000", 11278 => "0000000000000000", 11279 => "0000000000000000", 11280 => "0000000000000000", 11281 => "0000000000000000", 11282 => "0000000000000000", 11283 => "0000000000000000", 11284 => "0000000000000000", 11285 => "0000000000000000", 11286 => "0000000000000000", 11287 => "0000000000000000", 11288 => "0000000000000000", 11289 => "0000000000000000", 11290 => "0000000000000000", 11291 => "0000000000000000", 11292 => "0000000000000000", 11293 => "0000000000000000", 11294 => "0000000000000000", 11295 => "0000000000000000", 11296 => "0000000000000000", 11297 => "0000000000000000", 11298 => "0000000000000000", 11299 => "0000000000000000", 11300 => "0000000000000000", 11301 => "0000000000000000", 11302 => "0000000000000000", 11303 => "0000000000000000", 11304 => "0000000000000000", 11305 => "0000000000000000", 11306 => "0000000000000000", 11307 => "0000000000000000", 11308 => "0000000000000000", 11309 => "0000000000000000", 11310 => "0000000000000000", 11311 => "0000000000000000", 11312 => "0000000000000000", 11313 => "0000000000000000", 11314 => "0000000000000000", 11315 => "0000000000000000", 11316 => "0000000000000000", 11317 => "0000000000000000", 11318 => "0000000000000000", 11319 => "0000000000000000", 11320 => "0000000000000000", 11321 => "0000000000000000", 11322 => "0000000000000000", 11323 => "0000000000000000", 11324 => "0000000000000000", 11325 => "0000000000000000", 11326 => "0000000000000000", 11327 => "0000000000000000", 11328 => "0000000000000000", 11329 => "0000000000000000", 11330 => "0000000000000000", 11331 => "0000000000000000", 11332 => "0000000000000000", 11333 => "0000000000000000", 11334 => "0000000000000000", 11335 => "0000000000000000", 11336 => "0000000000000000", 11337 => "0000000000000000", 11338 => "0000000000000000", 11339 => "0000000000000000", 11340 => "0000000000000000", 11341 => "0000000000000000", 11342 => "0000000000000000", 11343 => "0000000000000000", 11344 => "0000000000000000", 11345 => "0000000000000000", 11346 => "0000000000000000", 11347 => "0000000000000000", 11348 => "0000000000000000", 11349 => "0000000000000000", 11350 => "0000000000000000", 11351 => "0000000000000000", 11352 => "0000000000000000", 11353 => "0000000000000000", 11354 => "0000000000000000", 11355 => "0000000000000000", 11356 => "0000000000000000", 11357 => "0000000000000000", 11358 => "0000000000000000", 11359 => "0000000000000000", 11360 => "0000000000000000", 11361 => "0000000000000000", 11362 => "0000000000000000", 11363 => "0000000000000000", 11364 => "0000000000000000", 11365 => "0000000000000000", 11366 => "0000000000000000", 11367 => "0000000000000000", 11368 => "0000000000000000", 11369 => "0000000000000000", 11370 => "0000000000000000", 11371 => "0000000000000000", 11372 => "0000000000000000", 11373 => "0000000000000000", 11374 => "0000000000000000", 11375 => "0000000000000000", 11376 => "0000000000000000", 11377 => "0000000000000000", 11378 => "0000000000000000", 11379 => "0000000000000000", 11380 => "0000000000000000", 11381 => "0000000000000000", 11382 => "0000000000000000", 11383 => "0000000000000000", 11384 => "0000000000000000", 11385 => "0000000000000000", 11386 => "0000000000000000", 11387 => "0000000000000000", 11388 => "0000000000000000", 11389 => "0000000000000000", 11390 => "0000000000000000", 11391 => "0000000000000000", 11392 => "0000000000000000", 11393 => "0000000000000000", 11394 => "0000000000000000", 11395 => "0000000000000000", 11396 => "0000000000000000", 11397 => "0000000000000000", 11398 => "0000000000000000", 11399 => "0000000000000000", 11400 => "0000000000000000", 11401 => "0000000000000000", 11402 => "0000000000000000", 11403 => "0000000000000000", 11404 => "0000000000000000", 11405 => "0000000000000000", 11406 => "0000000000000000", 11407 => "0000000000000000", 11408 => "0000000000000000", 11409 => "0000000000000000", 11410 => "0000000000000000", 11411 => "0000000000000000", 11412 => "0000000000000000", 11413 => "0000000000000000", 11414 => "0000000000000000", 11415 => "0000000000000000", 11416 => "0000000000000000", 11417 => "0000000000000000", 11418 => "0000000000000000", 11419 => "0000000000000000", 11420 => "0000000000000000", 11421 => "0000000000000000", 11422 => "0000000000000000", 11423 => "0000000000000000", 11424 => "0000000000000000", 11425 => "0000000000000000", 11426 => "0000000000000000", 11427 => "0000000000000000", 11428 => "0000000000000000", 11429 => "0000000000000000", 11430 => "0000000000000000", 11431 => "0000000000000000", 11432 => "0000000000000000", 11433 => "0000000000000000", 11434 => "0000000000000000", 11435 => "0000000000000000", 11436 => "0000000000000000", 11437 => "0000000000000000", 11438 => "0000000000000000", 11439 => "0000000000000000", 11440 => "0000000000000000", 11441 => "0000000000000000", 11442 => "0000000000000000", 11443 => "0000000000000000", 11444 => "0000000000000000", 11445 => "0000000000000000", 11446 => "0000000000000000", 11447 => "0000000000000000", 11448 => "0000000000000000", 11449 => "0000000000000000", 11450 => "0000000000000000", 11451 => "0000000000000000", 11452 => "0000000000000000", 11453 => "0000000000000000", 11454 => "0000000000000000", 11455 => "0000000000000000", 11456 => "0000000000000000", 11457 => "0000000000000000", 11458 => "0000000000000000", 11459 => "0000000000000000", 11460 => "0000000000000000", 11461 => "0000000000000000", 11462 => "0000000000000000", 11463 => "0000000000000000", 11464 => "0000000000000000", 11465 => "0000000000000000", 11466 => "0000000000000000", 11467 => "0000000000000000", 11468 => "0000000000000000", 11469 => "0000000000000000", 11470 => "0000000000000000", 11471 => "0000000000000000", 11472 => "0000000000000000", 11473 => "0000000000000000", 11474 => "0000000000000000", 11475 => "0000000000000000", 11476 => "0000000000000000", 11477 => "0000000000000000", 11478 => "0000000000000000", 11479 => "0000000000000000", 11480 => "0000000000000000", 11481 => "0000000000000000", 11482 => "0000000000000000", 11483 => "0000000000000000", 11484 => "0000000000000000", 11485 => "0000000000000000", 11486 => "0000000000000000", 11487 => "0000000000000000", 11488 => "0000000000000000", 11489 => "0000000000000000", 11490 => "0000000000000000", 11491 => "0000000000000000", 11492 => "0000000000000000", 11493 => "0000000000000000", 11494 => "0000000000000000", 11495 => "0000000000000000", 11496 => "0000000000000000", 11497 => "0000000000000000", 11498 => "0000000000000000", 11499 => "0000000000000000", 11500 => "0000000000000000", 11501 => "0000000000000000", 11502 => "0000000000000000", 11503 => "0000000000000000", 11504 => "0000000000000000", 11505 => "0000000000000000", 11506 => "0000000000000000", 11507 => "0000000000000000", 11508 => "0000000000000000", 11509 => "0000000000000000", 11510 => "0000000000000000", 11511 => "0000000000000000", 11512 => "0000000000000000", 11513 => "0000000000000000", 11514 => "0000000000000000", 11515 => "0000000000000000", 11516 => "0000000000000000", 11517 => "0000000000000000", 11518 => "0000000000000000", 11519 => "0000000000000000", 11520 => "0000000000000000", 11521 => "0000000000000000", 11522 => "0000000000000000", 11523 => "0000000000000000", 11524 => "0000000000000000", 11525 => "0000000000000000", 11526 => "0000000000000000", 11527 => "0000000000000000", 11528 => "0000000000000000", 11529 => "0000000000000000", 11530 => "0000000000000000", 11531 => "0000000000000000", 11532 => "0000000000000000", 11533 => "0000000000000000", 11534 => "0000000000000000", 11535 => "0000000000000000", 11536 => "0000000000000000", 11537 => "0000000000000000", 11538 => "0000000000000000", 11539 => "0000000000000000", 11540 => "0000000000000000", 11541 => "0000000000000000", 11542 => "0000000000000000", 11543 => "0000000000000000", 11544 => "0000000000000000", 11545 => "0000000000000000", 11546 => "0000000000000000", 11547 => "0000000000000000", 11548 => "0000000000000000", 11549 => "0000000000000000", 11550 => "0000000000000000", 11551 => "0000000000000000", 11552 => "0000000000000000", 11553 => "0000000000000000", 11554 => "0000000000000000", 11555 => "0000000000000000", 11556 => "0000000000000000", 11557 => "0000000000000000", 11558 => "0000000000000000", 11559 => "0000000000000000", 11560 => "0000000000000000", 11561 => "0000000000000000", 11562 => "0000000000000000", 11563 => "0000000000000000", 11564 => "0000000000000000", 11565 => "0000000000000000", 11566 => "0000000000000000", 11567 => "0000000000000000", 11568 => "0000000000000000", 11569 => "0000000000000000", 11570 => "0000000000000000", 11571 => "0000000000000000", 11572 => "0000000000000000", 11573 => "0000000000000000", 11574 => "0000000000000000", 11575 => "0000000000000000", 11576 => "0000000000000000", 11577 => "0000000000000000", 11578 => "0000000000000000", 11579 => "0000000000000000", 11580 => "0000000000000000", 11581 => "0000000000000000", 11582 => "0000000000000000", 11583 => "0000000000000000", 11584 => "0000000000000000", 11585 => "0000000000000000", 11586 => "0000000000000000", 11587 => "0000000000000000", 11588 => "0000000000000000", 11589 => "0000000000000000", 11590 => "0000000000000000", 11591 => "0000000000000000", 11592 => "0000000000000000", 11593 => "0000000000000000", 11594 => "0000000000000000", 11595 => "0000000000000000", 11596 => "0000000000000000", 11597 => "0000000000000000", 11598 => "0000000000000000", 11599 => "0000000000000000", 11600 => "0000000000000000", 11601 => "0000000000000000", 11602 => "0000000000000000", 11603 => "0000000000000000", 11604 => "0000000000000000", 11605 => "0000000000000000", 11606 => "0000000000000000", 11607 => "0000000000000000", 11608 => "0000000000000000", 11609 => "0000000000000000", 11610 => "0000000000000000", 11611 => "0000000000000000", 11612 => "0000000000000000", 11613 => "0000000000000000", 11614 => "0000000000000000", 11615 => "0000000000000000", 11616 => "0000000000000000", 11617 => "0000000000000000", 11618 => "0000000000000000", 11619 => "0000000000000000", 11620 => "0000000000000000", 11621 => "0000000000000000", 11622 => "0000000000000000", 11623 => "0000000000000000", 11624 => "0000000000000000", 11625 => "0000000000000000", 11626 => "0000000000000000", 11627 => "0000000000000000", 11628 => "0000000000000000", 11629 => "0000000000000000", 11630 => "0000000000000000", 11631 => "0000000000000000", 11632 => "0000000000000000", 11633 => "0000000000000000", 11634 => "0000000000000000", 11635 => "0000000000000000", 11636 => "0000000000000000", 11637 => "0000000000000000", 11638 => "0000000000000000", 11639 => "0000000000000000", 11640 => "0000000000000000", 11641 => "0000000000000000", 11642 => "0000000000000000", 11643 => "0000000000000000", 11644 => "0000000000000000", 11645 => "0000000000000000", 11646 => "0000000000000000", 11647 => "0000000000000000", 11648 => "0000000000000000", 11649 => "0000000000000000", 11650 => "0000000000000000", 11651 => "0000000000000000", 11652 => "0000000000000000", 11653 => "0000000000000000", 11654 => "0000000000000000", 11655 => "0000000000000000", 11656 => "0000000000000000", 11657 => "0000000000000000", 11658 => "0000000000000000", 11659 => "0000000000000000", 11660 => "0000000000000000", 11661 => "0000000000000000", 11662 => "0000000000000000", 11663 => "0000000000000000", 11664 => "0000000000000000", 11665 => "0000000000000000", 11666 => "0000000000000000", 11667 => "0000000000000000", 11668 => "0000000000000000", 11669 => "0000000000000000", 11670 => "0000000000000000", 11671 => "0000000000000000", 11672 => "0000000000000000", 11673 => "0000000000000000", 11674 => "0000000000000000", 11675 => "0000000000000000", 11676 => "0000000000000000", 11677 => "0000000000000000", 11678 => "0000000000000000", 11679 => "0000000000000000", 11680 => "0000000000000000", 11681 => "0000000000000000", 11682 => "0000000000000000", 11683 => "0000000000000000", 11684 => "0000000000000000", 11685 => "0000000000000000", 11686 => "0000000000000000", 11687 => "0000000000000000", 11688 => "0000000000000000", 11689 => "0000000000000000", 11690 => "0000000000000000", 11691 => "0000000000000000", 11692 => "0000000000000000", 11693 => "0000000000000000", 11694 => "0000000000000000", 11695 => "0000000000000000", 11696 => "0000000000000000", 11697 => "0000000000000000", 11698 => "0000000000000000", 11699 => "0000000000000000", 11700 => "0000000000000000", 11701 => "0000000000000000", 11702 => "0000000000000000", 11703 => "0000000000000000", 11704 => "0000000000000000", 11705 => "0000000000000000", 11706 => "0000000000000000", 11707 => "0000000000000000", 11708 => "0000000000000000", 11709 => "0000000000000000", 11710 => "0000000000000000", 11711 => "0000000000000000", 11712 => "0000000000000000", 11713 => "0000000000000000", 11714 => "0000000000000000", 11715 => "0000000000000000", 11716 => "0000000000000000", 11717 => "0000000000000000", 11718 => "0000000000000000", 11719 => "0000000000000000", 11720 => "0000000000000000", 11721 => "0000000000000000", 11722 => "0000000000000000", 11723 => "0000000000000000", 11724 => "0000000000000000", 11725 => "0000000000000000", 11726 => "0000000000000000", 11727 => "0000000000000000", 11728 => "0000000000000000", 11729 => "0000000000000000", 11730 => "0000000000000000", 11731 => "0000000000000000", 11732 => "0000000000000000", 11733 => "0000000000000000", 11734 => "0000000000000000", 11735 => "0000000000000000", 11736 => "0000000000000000", 11737 => "0000000000000000", 11738 => "0000000000000000", 11739 => "0000000000000000", 11740 => "0000000000000000", 11741 => "0000000000000000", 11742 => "0000000000000000", 11743 => "0000000000000000", 11744 => "0000000000000000", 11745 => "0000000000000000", 11746 => "0000000000000000", 11747 => "0000000000000000", 11748 => "0000000000000000", 11749 => "0000000000000000", 11750 => "0000000000000000", 11751 => "0000000000000000", 11752 => "0000000000000000", 11753 => "0000000000000000", 11754 => "0000000000000000", 11755 => "0000000000000000", 11756 => "0000000000000000", 11757 => "0000000000000000", 11758 => "0000000000000000", 11759 => "0000000000000000", 11760 => "0000000000000000", 11761 => "0000000000000000", 11762 => "0000000000000000", 11763 => "0000000000000000", 11764 => "0000000000000000", 11765 => "0000000000000000", 11766 => "0000000000000000", 11767 => "0000000000000000", 11768 => "0000000000000000", 11769 => "0000000000000000", 11770 => "0000000000000000", 11771 => "0000000000000000", 11772 => "0000000000000000", 11773 => "0000000000000000", 11774 => "0000000000000000", 11775 => "0000000000000000", 11776 => "0000000000000000", 11777 => "0000000000000000", 11778 => "0000000000000000", 11779 => "0000000000000000", 11780 => "0000000000000000", 11781 => "0000000000000000", 11782 => "0000000000000000", 11783 => "0000000000000000", 11784 => "0000000000000000", 11785 => "0000000000000000", 11786 => "0000000000000000", 11787 => "0000000000000000", 11788 => "0000000000000000", 11789 => "0000000000000000", 11790 => "0000000000000000", 11791 => "0000000000000000", 11792 => "0000000000000000", 11793 => "0000000000000000", 11794 => "0000000000000000", 11795 => "0000000000000000", 11796 => "0000000000000000", 11797 => "0000000000000000", 11798 => "0000000000000000", 11799 => "0000000000000000", 11800 => "0000000000000000", 11801 => "0000000000000000", 11802 => "0000000000000000", 11803 => "0000000000000000", 11804 => "0000000000000000", 11805 => "0000000000000000", 11806 => "0000000000000000", 11807 => "0000000000000000", 11808 => "0000000000000000", 11809 => "0000000000000000", 11810 => "0000000000000000", 11811 => "0000000000000000", 11812 => "0000000000000000", 11813 => "0000000000000000", 11814 => "0000000000000000", 11815 => "0000000000000000", 11816 => "0000000000000000", 11817 => "0000000000000000", 11818 => "0000000000000000", 11819 => "0000000000000000", 11820 => "0000000000000000", 11821 => "0000000000000000", 11822 => "0000000000000000", 11823 => "0000000000000000", 11824 => "0000000000000000", 11825 => "0000000000000000", 11826 => "0000000000000000", 11827 => "0000000000000000", 11828 => "0000000000000000", 11829 => "0000000000000000", 11830 => "0000000000000000", 11831 => "0000000000000000", 11832 => "0000000000000000", 11833 => "0000000000000000", 11834 => "0000000000000000", 11835 => "0000000000000000", 11836 => "0000000000000000", 11837 => "0000000000000000", 11838 => "0000000000000000", 11839 => "0000000000000000", 11840 => "0000000000000000", 11841 => "0000000000000000", 11842 => "0000000000000000", 11843 => "0000000000000000", 11844 => "0000000000000000", 11845 => "0000000000000000", 11846 => "0000000000000000", 11847 => "0000000000000000", 11848 => "0000000000000000", 11849 => "0000000000000000", 11850 => "0000000000000000", 11851 => "0000000000000000", 11852 => "0000000000000000", 11853 => "0000000000000000", 11854 => "0000000000000000", 11855 => "0000000000000000", 11856 => "0000000000000000", 11857 => "0000000000000000", 11858 => "0000000000000000", 11859 => "0000000000000000", 11860 => "0000000000000000", 11861 => "0000000000000000", 11862 => "0000000000000000", 11863 => "0000000000000000", 11864 => "0000000000000000", 11865 => "0000000000000000", 11866 => "0000000000000000", 11867 => "0000000000000000", 11868 => "0000000000000000", 11869 => "0000000000000000", 11870 => "0000000000000000", 11871 => "0000000000000000", 11872 => "0000000000000000", 11873 => "0000000000000000", 11874 => "0000000000000000", 11875 => "0000000000000000", 11876 => "0000000000000000", 11877 => "0000000000000000", 11878 => "0000000000000000", 11879 => "0000000000000000", 11880 => "0000000000000000", 11881 => "0000000000000000", 11882 => "0000000000000000", 11883 => "0000000000000000", 11884 => "0000000000000000", 11885 => "0000000000000000", 11886 => "0000000000000000", 11887 => "0000000000000000", 11888 => "0000000000000000", 11889 => "0000000000000000", 11890 => "0000000000000000", 11891 => "0000000000000000", 11892 => "0000000000000000", 11893 => "0000000000000000", 11894 => "0000000000000000", 11895 => "0000000000000000", 11896 => "0000000000000000", 11897 => "0000000000000000", 11898 => "0000000000000000", 11899 => "0000000000000000", 11900 => "0000000000000000", 11901 => "0000000000000000", 11902 => "0000000000000000", 11903 => "0000000000000000", 11904 => "0000000000000000", 11905 => "0000000000000000", 11906 => "0000000000000000", 11907 => "0000000000000000", 11908 => "0000000000000000", 11909 => "0000000000000000", 11910 => "0000000000000000", 11911 => "0000000000000000", 11912 => "0000000000000000", 11913 => "0000000000000000", 11914 => "0000000000000000", 11915 => "0000000000000000", 11916 => "0000000000000000", 11917 => "0000000000000000", 11918 => "0000000000000000", 11919 => "0000000000000000", 11920 => "0000000000000000", 11921 => "0000000000000000", 11922 => "0000000000000000", 11923 => "0000000000000000", 11924 => "0000000000000000", 11925 => "0000000000000000", 11926 => "0000000000000000", 11927 => "0000000000000000", 11928 => "0000000000000000", 11929 => "0000000000000000", 11930 => "0000000000000000", 11931 => "0000000000000000", 11932 => "0000000000000000", 11933 => "0000000000000000", 11934 => "0000000000000000", 11935 => "0000000000000000", 11936 => "0000000000000000", 11937 => "0000000000000000", 11938 => "0000000000000000", 11939 => "0000000000000000", 11940 => "0000000000000000", 11941 => "0000000000000000", 11942 => "0000000000000000", 11943 => "0000000000000000", 11944 => "0000000000000000", 11945 => "0000000000000000", 11946 => "0000000000000000", 11947 => "0000000000000000", 11948 => "0000000000000000", 11949 => "0000000000000000", 11950 => "0000000000000000", 11951 => "0000000000000000", 11952 => "0000000000000000", 11953 => "0000000000000000", 11954 => "0000000000000000", 11955 => "0000000000000000", 11956 => "0000000000000000", 11957 => "0000000000000000", 11958 => "0000000000000000", 11959 => "0000000000000000", 11960 => "0000000000000000", 11961 => "0000000000000000", 11962 => "0000000000000000", 11963 => "0000000000000000", 11964 => "0000000000000000", 11965 => "0000000000000000", 11966 => "0000000000000000", 11967 => "0000000000000000", 11968 => "0000000000000000", 11969 => "0000000000000000", 11970 => "0000000000000000", 11971 => "0000000000000000", 11972 => "0000000000000000", 11973 => "0000000000000000", 11974 => "0000000000000000", 11975 => "0000000000000000", 11976 => "0000000000000000", 11977 => "0000000000000000", 11978 => "0000000000000000", 11979 => "0000000000000000", 11980 => "0000000000000000", 11981 => "0000000000000000", 11982 => "0000000000000000", 11983 => "0000000000000000", 11984 => "0000000000000000", 11985 => "0000000000000000", 11986 => "0000000000000000", 11987 => "0000000000000000", 11988 => "0000000000000000", 11989 => "0000000000000000", 11990 => "0000000000000000", 11991 => "0000000000000000", 11992 => "0000000000000000", 11993 => "0000000000000000", 11994 => "0000000000000000", 11995 => "0000000000000000", 11996 => "0000000000000000", 11997 => "0000000000000000", 11998 => "0000000000000000", 11999 => "0000000000000000", 12000 => "0000000000000000", 12001 => "0000000000000000", 12002 => "0000000000000000", 12003 => "0000000000000000", 12004 => "0000000000000000", 12005 => "0000000000000000", 12006 => "0000000000000000", 12007 => "0000000000000000", 12008 => "0000000000000000", 12009 => "0000000000000000", 12010 => "0000000000000000", 12011 => "0000000000000000", 12012 => "0000000000000000", 12013 => "0000000000000000", 12014 => "0000000000000000", 12015 => "0000000000000000", 12016 => "0000000000000000", 12017 => "0000000000000000", 12018 => "0000000000000000", 12019 => "0000000000000000", 12020 => "0000000000000000", 12021 => "0000000000000000", 12022 => "0000000000000000", 12023 => "0000000000000000", 12024 => "0000000000000000", 12025 => "0000000000000000", 12026 => "0000000000000000", 12027 => "0000000000000000", 12028 => "0000000000000000", 12029 => "0000000000000000", 12030 => "0000000000000000", 12031 => "0000000000000000", 12032 => "0000000000000000", 12033 => "0000000000000000", 12034 => "0000000000000000", 12035 => "0000000000000000", 12036 => "0000000000000000", 12037 => "0000000000000000", 12038 => "0000000000000000", 12039 => "0000000000000000", 12040 => "0000000000000000", 12041 => "0000000000000000", 12042 => "0000000000000000", 12043 => "0000000000000000", 12044 => "0000000000000000", 12045 => "0000000000000000", 12046 => "0000000000000000", 12047 => "0000000000000000", 12048 => "0000000000000000", 12049 => "0000000000000000", 12050 => "0000000000000000", 12051 => "0000000000000000", 12052 => "0000000000000000", 12053 => "0000000000000000", 12054 => "0000000000000000", 12055 => "0000000000000000", 12056 => "0000000000000000", 12057 => "0000000000000000", 12058 => "0000000000000000", 12059 => "0000000000000000", 12060 => "0000000000000000", 12061 => "0000000000000000", 12062 => "0000000000000000", 12063 => "0000000000000000", 12064 => "0000000000000000", 12065 => "0000000000000000", 12066 => "0000000000000000", 12067 => "0000000000000000", 12068 => "0000000000000000", 12069 => "0000000000000000", 12070 => "0000000000000000", 12071 => "0000000000000000", 12072 => "0000000000000000", 12073 => "0000000000000000", 12074 => "0000000000000000", 12075 => "0000000000000000", 12076 => "0000000000000000", 12077 => "0000000000000000", 12078 => "0000000000000000", 12079 => "0000000000000000", 12080 => "0000000000000000", 12081 => "0000000000000000", 12082 => "0000000000000000", 12083 => "0000000000000000", 12084 => "0000000000000000", 12085 => "0000000000000000", 12086 => "0000000000000000", 12087 => "0000000000000000", 12088 => "0000000000000000", 12089 => "0000000000000000", 12090 => "0000000000000000", 12091 => "0000000000000000", 12092 => "0000000000000000", 12093 => "0000000000000000", 12094 => "0000000000000000", 12095 => "0000000000000000", 12096 => "0000000000000000", 12097 => "0000000000000000", 12098 => "0000000000000000", 12099 => "0000000000000000", 12100 => "0000000000000000", 12101 => "0000000000000000", 12102 => "0000000000000000", 12103 => "0000000000000000", 12104 => "0000000000000000", 12105 => "0000000000000000", 12106 => "0000000000000000", 12107 => "0000000000000000", 12108 => "0000000000000000", 12109 => "0000000000000000", 12110 => "0000000000000000", 12111 => "0000000000000000", 12112 => "0000000000000000", 12113 => "0000000000000000", 12114 => "0000000000000000", 12115 => "0000000000000000", 12116 => "0000000000000000", 12117 => "0000000000000000", 12118 => "0000000000000000", 12119 => "0000000000000000", 12120 => "0000000000000000", 12121 => "0000000000000000", 12122 => "0000000000000000", 12123 => "0000000000000000", 12124 => "0000000000000000", 12125 => "0000000000000000", 12126 => "0000000000000000", 12127 => "0000000000000000", 12128 => "0000000000000000", 12129 => "0000000000000000", 12130 => "0000000000000000", 12131 => "0000000000000000", 12132 => "0000000000000000", 12133 => "0000000000000000", 12134 => "0000000000000000", 12135 => "0000000000000000", 12136 => "0000000000000000", 12137 => "0000000000000000", 12138 => "0000000000000000", 12139 => "0000000000000000", 12140 => "0000000000000000", 12141 => "0000000000000000", 12142 => "0000000000000000", 12143 => "0000000000000000", 12144 => "0000000000000000", 12145 => "0000000000000000", 12146 => "0000000000000000", 12147 => "0000000000000000", 12148 => "0000000000000000", 12149 => "0000000000000000", 12150 => "0000000000000000", 12151 => "0000000000000000", 12152 => "0000000000000000", 12153 => "0000000000000000", 12154 => "0000000000000000", 12155 => "0000000000000000", 12156 => "0000000000000000", 12157 => "0000000000000000", 12158 => "0000000000000000", 12159 => "0000000000000000", 12160 => "0000000000000000", 12161 => "0000000000000000", 12162 => "0000000000000000", 12163 => "0000000000000000", 12164 => "0000000000000000", 12165 => "0000000000000000", 12166 => "0000000000000000", 12167 => "0000000000000000", 12168 => "0000000000000000", 12169 => "0000000000000000", 12170 => "0000000000000000", 12171 => "0000000000000000", 12172 => "0000000000000000", 12173 => "0000000000000000", 12174 => "0000000000000000", 12175 => "0000000000000000", 12176 => "0000000000000000", 12177 => "0000000000000000", 12178 => "0000000000000000", 12179 => "0000000000000000", 12180 => "0000000000000000", 12181 => "0000000000000000", 12182 => "0000000000000000", 12183 => "0000000000000000", 12184 => "0000000000000000", 12185 => "0000000000000000", 12186 => "0000000000000000", 12187 => "0000000000000000", 12188 => "0000000000000000", 12189 => "0000000000000000", 12190 => "0000000000000000", 12191 => "0000000000000000", 12192 => "0000000000000000", 12193 => "0000000000000000", 12194 => "0000000000000000", 12195 => "0000000000000000", 12196 => "0000000000000000", 12197 => "0000000000000000", 12198 => "0000000000000000", 12199 => "0000000000000000", 12200 => "0000000000000000", 12201 => "0000000000000000", 12202 => "0000000000000000", 12203 => "0000000000000000", 12204 => "0000000000000000", 12205 => "0000000000000000", 12206 => "0000000000000000", 12207 => "0000000000000000", 12208 => "0000000000000000", 12209 => "0000000000000000", 12210 => "0000000000000000", 12211 => "0000000000000000", 12212 => "0000000000000000", 12213 => "0000000000000000", 12214 => "0000000000000000", 12215 => "0000000000000000", 12216 => "0000000000000000", 12217 => "0000000000000000", 12218 => "0000000000000000", 12219 => "0000000000000000", 12220 => "0000000000000000", 12221 => "0000000000000000", 12222 => "0000000000000000", 12223 => "0000000000000000", 12224 => "0000000000000000", 12225 => "0000000000000000", 12226 => "0000000000000000", 12227 => "0000000000000000", 12228 => "0000000000000000", 12229 => "0000000000000000", 12230 => "0000000000000000", 12231 => "0000000000000000", 12232 => "0000000000000000", 12233 => "0000000000000000", 12234 => "0000000000000000", 12235 => "0000000000000000", 12236 => "0000000000000000", 12237 => "0000000000000000", 12238 => "0000000000000000", 12239 => "0000000000000000", 12240 => "0000000000000000", 12241 => "0000000000000000", 12242 => "0000000000000000", 12243 => "0000000000000000", 12244 => "0000000000000000", 12245 => "0000000000000000", 12246 => "0000000000000000", 12247 => "0000000000000000", 12248 => "0000000000000000", 12249 => "0000000000000000", 12250 => "0000000000000000", 12251 => "0000000000000000", 12252 => "0000000000000000", 12253 => "0000000000000000", 12254 => "0000000000000000", 12255 => "0000000000000000", 12256 => "0000000000000000", 12257 => "0000000000000000", 12258 => "0000000000000000", 12259 => "0000000000000000", 12260 => "0000000000000000", 12261 => "0000000000000000", 12262 => "0000000000000000", 12263 => "0000000000000000", 12264 => "0000000000000000", 12265 => "0000000000000000", 12266 => "0000000000000000", 12267 => "0000000000000000", 12268 => "0000000000000000", 12269 => "0000000000000000", 12270 => "0000000000000000", 12271 => "0000000000000000", 12272 => "0000000000000000", 12273 => "0000000000000000", 12274 => "0000000000000000", 12275 => "0000000000000000", 12276 => "0000000000000000", 12277 => "0000000000000000", 12278 => "0000000000000000", 12279 => "0000000000000000", 12280 => "0000000000000000", 12281 => "0000000000000000", 12282 => "0000000000000000", 12283 => "0000000000000000", 12284 => "0000000000000000", 12285 => "0000000000000000", 12286 => "0000000000000000", 12287 => "0000000000000000", 12288 => "0000000000000000", 12289 => "0000000000000000", 12290 => "0000000000000000", 12291 => "0000000000000000", 12292 => "0000000000000000", 12293 => "0000000000000000", 12294 => "0000000000000000", 12295 => "0000000000000000", 12296 => "0000000000000000", 12297 => "0000000000000000", 12298 => "0000000000000000", 12299 => "0000000000000000", 12300 => "0000000000000000", 12301 => "0000000000000000", 12302 => "0000000000000000", 12303 => "0000000000000000", 12304 => "0000000000000000", 12305 => "0000000000000000", 12306 => "0000000000000000", 12307 => "0000000000000000", 12308 => "0000000000000000", 12309 => "0000000000000000", 12310 => "0000000000000000", 12311 => "0000000000000000", 12312 => "0000000000000000", 12313 => "0000000000000000", 12314 => "0000000000000000", 12315 => "0000000000000000", 12316 => "0000000000000000", 12317 => "0000000000000000", 12318 => "0000000000000000", 12319 => "0000000000000000", 12320 => "0000000000000000", 12321 => "0000000000000000", 12322 => "0000000000000000", 12323 => "0000000000000000", 12324 => "0000000000000000", 12325 => "0000000000000000", 12326 => "0000000000000000", 12327 => "0000000000000000", 12328 => "0000000000000000", 12329 => "0000000000000000", 12330 => "0000000000000000", 12331 => "0000000000000000", 12332 => "0000000000000000", 12333 => "0000000000000000", 12334 => "0000000000000000", 12335 => "0000000000000000", 12336 => "0000000000000000", 12337 => "0000000000000000", 12338 => "0000000000000000", 12339 => "0000000000000000", 12340 => "0000000000000000", 12341 => "0000000000000000", 12342 => "0000000000000000", 12343 => "0000000000000000", 12344 => "0000000000000000", 12345 => "0000000000000000", 12346 => "0000000000000000", 12347 => "0000000000000000", 12348 => "0000000000000000", 12349 => "0000000000000000", 12350 => "0000000000000000", 12351 => "0000000000000000", 12352 => "0000000000000000", 12353 => "0000000000000000", 12354 => "0000000000000000", 12355 => "0000000000000000", 12356 => "0000000000000000", 12357 => "0000000000000000", 12358 => "0000000000000000", 12359 => "0000000000000000", 12360 => "0000000000000000", 12361 => "0000000000000000", 12362 => "0000000000000000", 12363 => "0000000000000000", 12364 => "0000000000000000", 12365 => "0000000000000000", 12366 => "0000000000000000", 12367 => "0000000000000000", 12368 => "0000000000000000", 12369 => "0000000000000000", 12370 => "0000000000000000", 12371 => "0000000000000000", 12372 => "0000000000000000", 12373 => "0000000000000000", 12374 => "0000000000000000", 12375 => "0000000000000000", 12376 => "0000000000000000", 12377 => "0000000000000000", 12378 => "0000000000000000", 12379 => "0000000000000000", 12380 => "0000000000000000", 12381 => "0000000000000000", 12382 => "0000000000000000", 12383 => "0000000000000000", 12384 => "0000000000000000", 12385 => "0000000000000000", 12386 => "0000000000000000", 12387 => "0000000000000000", 12388 => "0000000000000000", 12389 => "0000000000000000", 12390 => "0000000000000000", 12391 => "0000000000000000", 12392 => "0000000000000000", 12393 => "0000000000000000", 12394 => "0000000000000000", 12395 => "0000000000000000", 12396 => "0000000000000000", 12397 => "0000000000000000", 12398 => "0000000000000000", 12399 => "0000000000000000", 12400 => "0000000000000000", 12401 => "0000000000000000", 12402 => "0000000000000000", 12403 => "0000000000000000", 12404 => "0000000000000000", 12405 => "0000000000000000", 12406 => "0000000000000000", 12407 => "0000000000000000", 12408 => "0000000000000000", 12409 => "0000000000000000", 12410 => "0000000000000000", 12411 => "0000000000000000", 12412 => "0000000000000000", 12413 => "0000000000000000", 12414 => "0000000000000000", 12415 => "0000000000000000", 12416 => "0000000000000000", 12417 => "0000000000000000", 12418 => "0000000000000000", 12419 => "0000000000000000", 12420 => "0000000000000000", 12421 => "0000000000000000", 12422 => "0000000000000000", 12423 => "0000000000000000", 12424 => "0000000000000000", 12425 => "0000000000000000", 12426 => "0000000000000000", 12427 => "0000000000000000", 12428 => "0000000000000000", 12429 => "0000000000000000", 12430 => "0000000000000000", 12431 => "0000000000000000", 12432 => "0000000000000000", 12433 => "0000000000000000", 12434 => "0000000000000000", 12435 => "0000000000000000", 12436 => "0000000000000000", 12437 => "0000000000000000", 12438 => "0000000000000000", 12439 => "0000000000000000", 12440 => "0000000000000000", 12441 => "0000000000000000", 12442 => "0000000000000000", 12443 => "0000000000000000", 12444 => "0000000000000000", 12445 => "0000000000000000", 12446 => "0000000000000000", 12447 => "0000000000000000", 12448 => "0000000000000000", 12449 => "0000000000000000", 12450 => "0000000000000000", 12451 => "0000000000000000", 12452 => "0000000000000000", 12453 => "0000000000000000", 12454 => "0000000000000000", 12455 => "0000000000000000", 12456 => "0000000000000000", 12457 => "0000000000000000", 12458 => "0000000000000000", 12459 => "0000000000000000", 12460 => "0000000000000000", 12461 => "0000000000000000", 12462 => "0000000000000000", 12463 => "0000000000000000", 12464 => "0000000000000000", 12465 => "0000000000000000", 12466 => "0000000000000000", 12467 => "0000000000000000", 12468 => "0000000000000000", 12469 => "0000000000000000", 12470 => "0000000000000000", 12471 => "0000000000000000", 12472 => "0000000000000000", 12473 => "0000000000000000", 12474 => "0000000000000000", 12475 => "0000000000000000", 12476 => "0000000000000000", 12477 => "0000000000000000", 12478 => "0000000000000000", 12479 => "0000000000000000", 12480 => "0000000000000000", 12481 => "0000000000000000", 12482 => "0000000000000000", 12483 => "0000000000000000", 12484 => "0000000000000000", 12485 => "0000000000000000", 12486 => "0000000000000000", 12487 => "0000000000000000", 12488 => "0000000000000000", 12489 => "0000000000000000", 12490 => "0000000000000000", 12491 => "0000000000000000", 12492 => "0000000000000000", 12493 => "0000000000000000", 12494 => "0000000000000000", 12495 => "0000000000000000", 12496 => "0000000000000000", 12497 => "0000000000000000", 12498 => "0000000000000000", 12499 => "0000000000000000", 12500 => "0000000000000000", 12501 => "0000000000000000", 12502 => "0000000000000000", 12503 => "0000000000000000", 12504 => "0000000000000000", 12505 => "0000000000000000", 12506 => "0000000000000000", 12507 => "0000000000000000", 12508 => "0000000000000000", 12509 => "0000000000000000", 12510 => "0000000000000000", 12511 => "0000000000000000", 12512 => "0000000000000000", 12513 => "0000000000000000", 12514 => "0000000000000000", 12515 => "0000000000000000", 12516 => "0000000000000000", 12517 => "0000000000000000", 12518 => "0000000000000000", 12519 => "0000000000000000", 12520 => "0000000000000000", 12521 => "0000000000000000", 12522 => "0000000000000000", 12523 => "0000000000000000", 12524 => "0000000000000000", 12525 => "0000000000000000", 12526 => "0000000000000000", 12527 => "0000000000000000", 12528 => "0000000000000000", 12529 => "0000000000000000", 12530 => "0000000000000000", 12531 => "0000000000000000", 12532 => "0000000000000000", 12533 => "0000000000000000", 12534 => "0000000000000000", 12535 => "0000000000000000", 12536 => "0000000000000000", 12537 => "0000000000000000", 12538 => "0000000000000000", 12539 => "0000000000000000", 12540 => "0000000000000000", 12541 => "0000000000000000", 12542 => "0000000000000000", 12543 => "0000000000000000", 12544 => "0000000000000000", 12545 => "0000000000000000", 12546 => "0000000000000000", 12547 => "0000000000000000", 12548 => "0000000000000000", 12549 => "0000000000000000", 12550 => "0000000000000000", 12551 => "0000000000000000", 12552 => "0000000000000000", 12553 => "0000000000000000", 12554 => "0000000000000000", 12555 => "0000000000000000", 12556 => "0000000000000000", 12557 => "0000000000000000", 12558 => "0000000000000000", 12559 => "0000000000000000", 12560 => "0000000000000000", 12561 => "0000000000000000", 12562 => "0000000000000000", 12563 => "0000000000000000", 12564 => "0000000000000000", 12565 => "0000000000000000", 12566 => "0000000000000000", 12567 => "0000000000000000", 12568 => "0000000000000000", 12569 => "0000000000000000", 12570 => "0000000000000000", 12571 => "0000000000000000", 12572 => "0000000000000000", 12573 => "0000000000000000", 12574 => "0000000000000000", 12575 => "0000000000000000", 12576 => "0000000000000000", 12577 => "0000000000000000", 12578 => "0000000000000000", 12579 => "0000000000000000", 12580 => "0000000000000000", 12581 => "0000000000000000", 12582 => "0000000000000000", 12583 => "0000000000000000", 12584 => "0000000000000000", 12585 => "0000000000000000", 12586 => "0000000000000000", 12587 => "0000000000000000", 12588 => "0000000000000000", 12589 => "0000000000000000", 12590 => "0000000000000000", 12591 => "0000000000000000", 12592 => "0000000000000000", 12593 => "0000000000000000", 12594 => "0000000000000000", 12595 => "0000000000000000", 12596 => "0000000000000000", 12597 => "0000000000000000", 12598 => "0000000000000000", 12599 => "0000000000000000", 12600 => "0000000000000000", 12601 => "0000000000000000", 12602 => "0000000000000000", 12603 => "0000000000000000", 12604 => "0000000000000000", 12605 => "0000000000000000", 12606 => "0000000000000000", 12607 => "0000000000000000", 12608 => "0000000000000000", 12609 => "0000000000000000", 12610 => "0000000000000000", 12611 => "0000000000000000", 12612 => "0000000000000000", 12613 => "0000000000000000", 12614 => "0000000000000000", 12615 => "0000000000000000", 12616 => "0000000000000000", 12617 => "0000000000000000", 12618 => "0000000000000000", 12619 => "0000000000000000", 12620 => "0000000000000000", 12621 => "0000000000000000", 12622 => "0000000000000000", 12623 => "0000000000000000", 12624 => "0000000000000000", 12625 => "0000000000000000", 12626 => "0000000000000000", 12627 => "0000000000000000", 12628 => "0000000000000000", 12629 => "0000000000000000", 12630 => "0000000000000000", 12631 => "0000000000000000", 12632 => "0000000000000000", 12633 => "0000000000000000", 12634 => "0000000000000000", 12635 => "0000000000000000", 12636 => "0000000000000000", 12637 => "0000000000000000", 12638 => "0000000000000000", 12639 => "0000000000000000", 12640 => "0000000000000000", 12641 => "0000000000000000", 12642 => "0000000000000000", 12643 => "0000000000000000", 12644 => "0000000000000000", 12645 => "0000000000000000", 12646 => "0000000000000000", 12647 => "0000000000000000", 12648 => "0000000000000000", 12649 => "0000000000000000", 12650 => "0000000000000000", 12651 => "0000000000000000", 12652 => "0000000000000000", 12653 => "0000000000000000", 12654 => "0000000000000000", 12655 => "0000000000000000", 12656 => "0000000000000000", 12657 => "0000000000000000", 12658 => "0000000000000000", 12659 => "0000000000000000", 12660 => "0000000000000000", 12661 => "0000000000000000", 12662 => "0000000000000000", 12663 => "0000000000000000", 12664 => "0000000000000000", 12665 => "0000000000000000", 12666 => "0000000000000000", 12667 => "0000000000000000", 12668 => "0000000000000000", 12669 => "0000000000000000", 12670 => "0000000000000000", 12671 => "0000000000000000", 12672 => "0000000000000000", 12673 => "0000000000000000", 12674 => "0000000000000000", 12675 => "0000000000000000", 12676 => "0000000000000000", 12677 => "0000000000000000", 12678 => "0000000000000000", 12679 => "0000000000000000", 12680 => "0000000000000000", 12681 => "0000000000000000", 12682 => "0000000000000000", 12683 => "0000000000000000", 12684 => "0000000000000000", 12685 => "0000000000000000", 12686 => "0000000000000000", 12687 => "0000000000000000", 12688 => "0000000000000000", 12689 => "0000000000000000", 12690 => "0000000000000000", 12691 => "0000000000000000", 12692 => "0000000000000000", 12693 => "0000000000000000", 12694 => "0000000000000000", 12695 => "0000000000000000", 12696 => "0000000000000000", 12697 => "0000000000000000", 12698 => "0000000000000000", 12699 => "0000000000000000", 12700 => "0000000000000000", 12701 => "0000000000000000", 12702 => "0000000000000000", 12703 => "0000000000000000", 12704 => "0000000000000000", 12705 => "0000000000000000", 12706 => "0000000000000000", 12707 => "0000000000000000", 12708 => "0000000000000000", 12709 => "0000000000000000", 12710 => "0000000000000000", 12711 => "0000000000000000", 12712 => "0000000000000000", 12713 => "0000000000000000", 12714 => "0000000000000000", 12715 => "0000000000000000", 12716 => "0000000000000000", 12717 => "0000000000000000", 12718 => "0000000000000000", 12719 => "0000000000000000", 12720 => "0000000000000000", 12721 => "0000000000000000", 12722 => "0000000000000000", 12723 => "0000000000000000", 12724 => "0000000000000000", 12725 => "0000000000000000", 12726 => "0000000000000000", 12727 => "0000000000000000", 12728 => "0000000000000000", 12729 => "0000000000000000", 12730 => "0000000000000000", 12731 => "0000000000000000", 12732 => "0000000000000000", 12733 => "0000000000000000", 12734 => "0000000000000000", 12735 => "0000000000000000", 12736 => "0000000000000000", 12737 => "0000000000000000", 12738 => "0000000000000000", 12739 => "0000000000000000", 12740 => "0000000000000000", 12741 => "0000000000000000", 12742 => "0000000000000000", 12743 => "0000000000000000", 12744 => "0000000000000000", 12745 => "0000000000000000", 12746 => "0000000000000000", 12747 => "0000000000000000", 12748 => "0000000000000000", 12749 => "0000000000000000", 12750 => "0000000000000000", 12751 => "0000000000000000", 12752 => "0000000000000000", 12753 => "0000000000000000", 12754 => "0000000000000000", 12755 => "0000000000000000", 12756 => "0000000000000000", 12757 => "0000000000000000", 12758 => "0000000000000000", 12759 => "0000000000000000", 12760 => "0000000000000000", 12761 => "0000000000000000", 12762 => "0000000000000000", 12763 => "0000000000000000", 12764 => "0000000000000000", 12765 => "0000000000000000", 12766 => "0000000000000000", 12767 => "0000000000000000", 12768 => "0000000000000000", 12769 => "0000000000000000", 12770 => "0000000000000000", 12771 => "0000000000000000", 12772 => "0000000000000000", 12773 => "0000000000000000", 12774 => "0000000000000000", 12775 => "0000000000000000", 12776 => "0000000000000000", 12777 => "0000000000000000", 12778 => "0000000000000000", 12779 => "0000000000000000", 12780 => "0000000000000000", 12781 => "0000000000000000", 12782 => "0000000000000000", 12783 => "0000000000000000", 12784 => "0000000000000000", 12785 => "0000000000000000", 12786 => "0000000000000000", 12787 => "0000000000000000", 12788 => "0000000000000000", 12789 => "0000000000000000", 12790 => "0000000000000000", 12791 => "0000000000000000", 12792 => "0000000000000000", 12793 => "0000000000000000", 12794 => "0000000000000000", 12795 => "0000000000000000", 12796 => "0000000000000000", 12797 => "0000000000000000", 12798 => "0000000000000000", 12799 => "0000000000000000", 12800 => "0000000000000000", 12801 => "0000000000000000", 12802 => "0000000000000000", 12803 => "0000000000000000", 12804 => "0000000000000000", 12805 => "0000000000000000", 12806 => "0000000000000000", 12807 => "0000000000000000", 12808 => "0000000000000000", 12809 => "0000000000000000", 12810 => "0000000000000000", 12811 => "0000000000000000", 12812 => "0000000000000000", 12813 => "0000000000000000", 12814 => "0000000000000000", 12815 => "0000000000000000", 12816 => "0000000000000000", 12817 => "0000000000000000", 12818 => "0000000000000000", 12819 => "0000000000000000", 12820 => "0000000000000000", 12821 => "0000000000000000", 12822 => "0000000000000000", 12823 => "0000000000000000", 12824 => "0000000000000000", 12825 => "0000000000000000", 12826 => "0000000000000000", 12827 => "0000000000000000", 12828 => "0000000000000000", 12829 => "0000000000000000", 12830 => "0000000000000000", 12831 => "0000000000000000", 12832 => "0000000000000000", 12833 => "0000000000000000", 12834 => "0000000000000000", 12835 => "0000000000000000", 12836 => "0000000000000000", 12837 => "0000000000000000", 12838 => "0000000000000000", 12839 => "0000000000000000", 12840 => "0000000000000000", 12841 => "0000000000000000", 12842 => "0000000000000000", 12843 => "0000000000000000", 12844 => "0000000000000000", 12845 => "0000000000000000", 12846 => "0000000000000000", 12847 => "0000000000000000", 12848 => "0000000000000000", 12849 => "0000000000000000", 12850 => "0000000000000000", 12851 => "0000000000000000", 12852 => "0000000000000000", 12853 => "0000000000000000", 12854 => "0000000000000000", 12855 => "0000000000000000", 12856 => "0000000000000000", 12857 => "0000000000000000", 12858 => "0000000000000000", 12859 => "0000000000000000", 12860 => "0000000000000000", 12861 => "0000000000000000", 12862 => "0000000000000000", 12863 => "0000000000000000", 12864 => "0000000000000000", 12865 => "0000000000000000", 12866 => "0000000000000000", 12867 => "0000000000000000", 12868 => "0000000000000000", 12869 => "0000000000000000", 12870 => "0000000000000000", 12871 => "0000000000000000", 12872 => "0000000000000000", 12873 => "0000000000000000", 12874 => "0000000000000000", 12875 => "0000000000000000", 12876 => "0000000000000000", 12877 => "0000000000000000", 12878 => "0000000000000000", 12879 => "0000000000000000", 12880 => "0000000000000000", 12881 => "0000000000000000", 12882 => "0000000000000000", 12883 => "0000000000000000", 12884 => "0000000000000000", 12885 => "0000000000000000", 12886 => "0000000000000000", 12887 => "0000000000000000", 12888 => "0000000000000000", 12889 => "0000000000000000", 12890 => "0000000000000000", 12891 => "0000000000000000", 12892 => "0000000000000000", 12893 => "0000000000000000", 12894 => "0000000000000000", 12895 => "0000000000000000", 12896 => "0000000000000000", 12897 => "0000000000000000", 12898 => "0000000000000000", 12899 => "0000000000000000", 12900 => "0000000000000000", 12901 => "0000000000000000", 12902 => "0000000000000000", 12903 => "0000000000000000", 12904 => "0000000000000000", 12905 => "0000000000000000", 12906 => "0000000000000000", 12907 => "0000000000000000", 12908 => "0000000000000000", 12909 => "0000000000000000", 12910 => "0000000000000000", 12911 => "0000000000000000", 12912 => "0000000000000000", 12913 => "0000000000000000", 12914 => "0000000000000000", 12915 => "0000000000000000", 12916 => "0000000000000000", 12917 => "0000000000000000", 12918 => "0000000000000000", 12919 => "0000000000000000", 12920 => "0000000000000000", 12921 => "0000000000000000", 12922 => "0000000000000000", 12923 => "0000000000000000", 12924 => "0000000000000000", 12925 => "0000000000000000", 12926 => "0000000000000000", 12927 => "0000000000000000", 12928 => "0000000000000000", 12929 => "0000000000000000", 12930 => "0000000000000000", 12931 => "0000000000000000", 12932 => "0000000000000000", 12933 => "0000000000000000", 12934 => "0000000000000000", 12935 => "0000000000000000", 12936 => "0000000000000000", 12937 => "0000000000000000", 12938 => "0000000000000000", 12939 => "0000000000000000", 12940 => "0000000000000000", 12941 => "0000000000000000", 12942 => "0000000000000000", 12943 => "0000000000000000", 12944 => "0000000000000000", 12945 => "0000000000000000", 12946 => "0000000000000000", 12947 => "0000000000000000", 12948 => "0000000000000000", 12949 => "0000000000000000", 12950 => "0000000000000000", 12951 => "0000000000000000", 12952 => "0000000000000000", 12953 => "0000000000000000", 12954 => "0000000000000000", 12955 => "0000000000000000", 12956 => "0000000000000000", 12957 => "0000000000000000", 12958 => "0000000000000000", 12959 => "0000000000000000", 12960 => "0000000000000000", 12961 => "0000000000000000", 12962 => "0000000000000000", 12963 => "0000000000000000", 12964 => "0000000000000000", 12965 => "0000000000000000", 12966 => "0000000000000000", 12967 => "0000000000000000", 12968 => "0000000000000000", 12969 => "0000000000000000", 12970 => "0000000000000000", 12971 => "0000000000000000", 12972 => "0000000000000000", 12973 => "0000000000000000", 12974 => "0000000000000000", 12975 => "0000000000000000", 12976 => "0000000000000000", 12977 => "0000000000000000", 12978 => "0000000000000000", 12979 => "0000000000000000", 12980 => "0000000000000000", 12981 => "0000000000000000", 12982 => "0000000000000000", 12983 => "0000000000000000", 12984 => "0000000000000000", 12985 => "0000000000000000", 12986 => "0000000000000000", 12987 => "0000000000000000", 12988 => "0000000000000000", 12989 => "0000000000000000", 12990 => "0000000000000000", 12991 => "0000000000000000", 12992 => "0000000000000000", 12993 => "0000000000000000", 12994 => "0000000000000000", 12995 => "0000000000000000", 12996 => "0000000000000000", 12997 => "0000000000000000", 12998 => "0000000000000000", 12999 => "0000000000000000", 13000 => "0000000000000000", 13001 => "0000000000000000", 13002 => "0000000000000000", 13003 => "0000000000000000", 13004 => "0000000000000000", 13005 => "0000000000000000", 13006 => "0000000000000000", 13007 => "0000000000000000", 13008 => "0000000000000000", 13009 => "0000000000000000", 13010 => "0000000000000000", 13011 => "0000000000000000", 13012 => "0000000000000000", 13013 => "0000000000000000", 13014 => "0000000000000000", 13015 => "0000000000000000", 13016 => "0000000000000000", 13017 => "0000000000000000", 13018 => "0000000000000000", 13019 => "0000000000000000", 13020 => "0000000000000000", 13021 => "0000000000000000", 13022 => "0000000000000000", 13023 => "0000000000000000", 13024 => "0000000000000000", 13025 => "0000000000000000", 13026 => "0000000000000000", 13027 => "0000000000000000", 13028 => "0000000000000000", 13029 => "0000000000000000", 13030 => "0000000000000000", 13031 => "0000000000000000", 13032 => "0000000000000000", 13033 => "0000000000000000", 13034 => "0000000000000000", 13035 => "0000000000000000", 13036 => "0000000000000000", 13037 => "0000000000000000", 13038 => "0000000000000000", 13039 => "0000000000000000", 13040 => "0000000000000000", 13041 => "0000000000000000", 13042 => "0000000000000000", 13043 => "0000000000000000", 13044 => "0000000000000000", 13045 => "0000000000000000", 13046 => "0000000000000000", 13047 => "0000000000000000", 13048 => "0000000000000000", 13049 => "0000000000000000", 13050 => "0000000000000000", 13051 => "0000000000000000", 13052 => "0000000000000000", 13053 => "0000000000000000", 13054 => "0000000000000000", 13055 => "0000000000000000", 13056 => "0000000000000000", 13057 => "0000000000000000", 13058 => "0000000000000000", 13059 => "0000000000000000", 13060 => "0000000000000000", 13061 => "0000000000000000", 13062 => "0000000000000000", 13063 => "0000000000000000", 13064 => "0000000000000000", 13065 => "0000000000000000", 13066 => "0000000000000000", 13067 => "0000000000000000", 13068 => "0000000000000000", 13069 => "0000000000000000", 13070 => "0000000000000000", 13071 => "0000000000000000", 13072 => "0000000000000000", 13073 => "0000000000000000", 13074 => "0000000000000000", 13075 => "0000000000000000", 13076 => "0000000000000000", 13077 => "0000000000000000", 13078 => "0000000000000000", 13079 => "0000000000000000", 13080 => "0000000000000000", 13081 => "0000000000000000", 13082 => "0000000000000000", 13083 => "0000000000000000", 13084 => "0000000000000000", 13085 => "0000000000000000", 13086 => "0000000000000000", 13087 => "0000000000000000", 13088 => "0000000000000000", 13089 => "0000000000000000", 13090 => "0000000000000000", 13091 => "0000000000000000", 13092 => "0000000000000000", 13093 => "0000000000000000", 13094 => "0000000000000000", 13095 => "0000000000000000", 13096 => "0000000000000000", 13097 => "0000000000000000", 13098 => "0000000000000000", 13099 => "0000000000000000", 13100 => "0000000000000000", 13101 => "0000000000000000", 13102 => "0000000000000000", 13103 => "0000000000000000", 13104 => "0000000000000000", 13105 => "0000000000000000", 13106 => "0000000000000000", 13107 => "0000000000000000", 13108 => "0000000000000000", 13109 => "0000000000000000", 13110 => "0000000000000000", 13111 => "0000000000000000", 13112 => "0000000000000000", 13113 => "0000000000000000", 13114 => "0000000000000000", 13115 => "0000000000000000", 13116 => "0000000000000000", 13117 => "0000000000000000", 13118 => "0000000000000000", 13119 => "0000000000000000", 13120 => "0000000000000000", 13121 => "0000000000000000", 13122 => "0000000000000000", 13123 => "0000000000000000", 13124 => "0000000000000000", 13125 => "0000000000000000", 13126 => "0000000000000000", 13127 => "0000000000000000", 13128 => "0000000000000000", 13129 => "0000000000000000", 13130 => "0000000000000000", 13131 => "0000000000000000", 13132 => "0000000000000000", 13133 => "0000000000000000", 13134 => "0000000000000000", 13135 => "0000000000000000", 13136 => "0000000000000000", 13137 => "0000000000000000", 13138 => "0000000000000000", 13139 => "0000000000000000", 13140 => "0000000000000000", 13141 => "0000000000000000", 13142 => "0000000000000000", 13143 => "0000000000000000", 13144 => "0000000000000000", 13145 => "0000000000000000", 13146 => "0000000000000000", 13147 => "0000000000000000", 13148 => "0000000000000000", 13149 => "0000000000000000", 13150 => "0000000000000000", 13151 => "0000000000000000", 13152 => "0000000000000000", 13153 => "0000000000000000", 13154 => "0000000000000000", 13155 => "0000000000000000", 13156 => "0000000000000000", 13157 => "0000000000000000", 13158 => "0000000000000000", 13159 => "0000000000000000", 13160 => "0000000000000000", 13161 => "0000000000000000", 13162 => "0000000000000000", 13163 => "0000000000000000", 13164 => "0000000000000000", 13165 => "0000000000000000", 13166 => "0000000000000000", 13167 => "0000000000000000", 13168 => "0000000000000000", 13169 => "0000000000000000", 13170 => "0000000000000000", 13171 => "0000000000000000", 13172 => "0000000000000000", 13173 => "0000000000000000", 13174 => "0000000000000000", 13175 => "0000000000000000", 13176 => "0000000000000000", 13177 => "0000000000000000", 13178 => "0000000000000000", 13179 => "0000000000000000", 13180 => "0000000000000000", 13181 => "0000000000000000", 13182 => "0000000000000000", 13183 => "0000000000000000", 13184 => "0000000000000000", 13185 => "0000000000000000", 13186 => "0000000000000000", 13187 => "0000000000000000", 13188 => "0000000000000000", 13189 => "0000000000000000", 13190 => "0000000000000000", 13191 => "0000000000000000", 13192 => "0000000000000000", 13193 => "0000000000000000", 13194 => "0000000000000000", 13195 => "0000000000000000", 13196 => "0000000000000000", 13197 => "0000000000000000", 13198 => "0000000000000000", 13199 => "0000000000000000", 13200 => "0000000000000000", 13201 => "0000000000000000", 13202 => "0000000000000000", 13203 => "0000000000000000", 13204 => "0000000000000000", 13205 => "0000000000000000", 13206 => "0000000000000000", 13207 => "0000000000000000", 13208 => "0000000000000000", 13209 => "0000000000000000", 13210 => "0000000000000000", 13211 => "0000000000000000", 13212 => "0000000000000000", 13213 => "0000000000000000", 13214 => "0000000000000000", 13215 => "0000000000000000", 13216 => "0000000000000000", 13217 => "0000000000000000", 13218 => "0000000000000000", 13219 => "0000000000000000", 13220 => "0000000000000000", 13221 => "0000000000000000", 13222 => "0000000000000000", 13223 => "0000000000000000", 13224 => "0000000000000000", 13225 => "0000000000000000", 13226 => "0000000000000000", 13227 => "0000000000000000", 13228 => "0000000000000000", 13229 => "0000000000000000", 13230 => "0000000000000000", 13231 => "0000000000000000", 13232 => "0000000000000000", 13233 => "0000000000000000", 13234 => "0000000000000000", 13235 => "0000000000000000", 13236 => "0000000000000000", 13237 => "0000000000000000", 13238 => "0000000000000000", 13239 => "0000000000000000", 13240 => "0000000000000000", 13241 => "0000000000000000", 13242 => "0000000000000000", 13243 => "0000000000000000", 13244 => "0000000000000000", 13245 => "0000000000000000", 13246 => "0000000000000000", 13247 => "0000000000000000", 13248 => "0000000000000000", 13249 => "0000000000000000", 13250 => "0000000000000000", 13251 => "0000000000000000", 13252 => "0000000000000000", 13253 => "0000000000000000", 13254 => "0000000000000000", 13255 => "0000000000000000", 13256 => "0000000000000000", 13257 => "0000000000000000", 13258 => "0000000000000000", 13259 => "0000000000000000", 13260 => "0000000000000000", 13261 => "0000000000000000", 13262 => "0000000000000000", 13263 => "0000000000000000", 13264 => "0000000000000000", 13265 => "0000000000000000", 13266 => "0000000000000000", 13267 => "0000000000000000", 13268 => "0000000000000000", 13269 => "0000000000000000", 13270 => "0000000000000000", 13271 => "0000000000000000", 13272 => "0000000000000000", 13273 => "0000000000000000", 13274 => "0000000000000000", 13275 => "0000000000000000", 13276 => "0000000000000000", 13277 => "0000000000000000", 13278 => "0000000000000000", 13279 => "0000000000000000", 13280 => "0000000000000000", 13281 => "0000000000000000", 13282 => "0000000000000000", 13283 => "0000000000000000", 13284 => "0000000000000000", 13285 => "0000000000000000", 13286 => "0000000000000000", 13287 => "0000000000000000", 13288 => "0000000000000000", 13289 => "0000000000000000", 13290 => "0000000000000000", 13291 => "0000000000000000", 13292 => "0000000000000000", 13293 => "0000000000000000", 13294 => "0000000000000000", 13295 => "0000000000000000", 13296 => "0000000000000000", 13297 => "0000000000000000", 13298 => "0000000000000000", 13299 => "0000000000000000", 13300 => "0000000000000000", 13301 => "0000000000000000", 13302 => "0000000000000000", 13303 => "0000000000000000", 13304 => "0000000000000000", 13305 => "0000000000000000", 13306 => "0000000000000000", 13307 => "0000000000000000", 13308 => "0000000000000000", 13309 => "0000000000000000", 13310 => "0000000000000000", 13311 => "0000000000000000", 13312 => "0000000000000000", 13313 => "0000000000000000", 13314 => "0000000000000000", 13315 => "0000000000000000", 13316 => "0000000000000000", 13317 => "0000000000000000", 13318 => "0000000000000000", 13319 => "0000000000000000", 13320 => "0000000000000000", 13321 => "0000000000000000", 13322 => "0000000000000000", 13323 => "0000000000000000", 13324 => "0000000000000000", 13325 => "0000000000000000", 13326 => "0000000000000000", 13327 => "0000000000000000", 13328 => "0000000000000000", 13329 => "0000000000000000", 13330 => "0000000000000000", 13331 => "0000000000000000", 13332 => "0000000000000000", 13333 => "0000000000000000", 13334 => "0000000000000000", 13335 => "0000000000000000", 13336 => "0000000000000000", 13337 => "0000000000000000", 13338 => "0000000000000000", 13339 => "0000000000000000", 13340 => "0000000000000000", 13341 => "0000000000000000", 13342 => "0000000000000000", 13343 => "0000000000000000", 13344 => "0000000000000000", 13345 => "0000000000000000", 13346 => "0000000000000000", 13347 => "0000000000000000", 13348 => "0000000000000000", 13349 => "0000000000000000", 13350 => "0000000000000000", 13351 => "0000000000000000", 13352 => "0000000000000000", 13353 => "0000000000000000", 13354 => "0000000000000000", 13355 => "0000000000000000", 13356 => "0000000000000000", 13357 => "0000000000000000", 13358 => "0000000000000000", 13359 => "0000000000000000", 13360 => "0000000000000000", 13361 => "0000000000000000", 13362 => "0000000000000000", 13363 => "0000000000000000", 13364 => "0000000000000000", 13365 => "0000000000000000", 13366 => "0000000000000000", 13367 => "0000000000000000", 13368 => "0000000000000000", 13369 => "0000000000000000", 13370 => "0000000000000000", 13371 => "0000000000000000", 13372 => "0000000000000000", 13373 => "0000000000000000", 13374 => "0000000000000000", 13375 => "0000000000000000", 13376 => "0000000000000000", 13377 => "0000000000000000", 13378 => "0000000000000000", 13379 => "0000000000000000", 13380 => "0000000000000000", 13381 => "0000000000000000", 13382 => "0000000000000000", 13383 => "0000000000000000", 13384 => "0000000000000000", 13385 => "0000000000000000", 13386 => "0000000000000000", 13387 => "0000000000000000", 13388 => "0000000000000000", 13389 => "0000000000000000", 13390 => "0000000000000000", 13391 => "0000000000000000", 13392 => "0000000000000000", 13393 => "0000000000000000", 13394 => "0000000000000000", 13395 => "0000000000000000", 13396 => "0000000000000000", 13397 => "0000000000000000", 13398 => "0000000000000000", 13399 => "0000000000000000", 13400 => "0000000000000000", 13401 => "0000000000000000", 13402 => "0000000000000000", 13403 => "0000000000000000", 13404 => "0000000000000000", 13405 => "0000000000000000", 13406 => "0000000000000000", 13407 => "0000000000000000", 13408 => "0000000000000000", 13409 => "0000000000000000", 13410 => "0000000000000000", 13411 => "0000000000000000", 13412 => "0000000000000000", 13413 => "0000000000000000", 13414 => "0000000000000000", 13415 => "0000000000000000", 13416 => "0000000000000000", 13417 => "0000000000000000", 13418 => "0000000000000000", 13419 => "0000000000000000", 13420 => "0000000000000000", 13421 => "0000000000000000", 13422 => "0000000000000000", 13423 => "0000000000000000", 13424 => "0000000000000000", 13425 => "0000000000000000", 13426 => "0000000000000000", 13427 => "0000000000000000", 13428 => "0000000000000000", 13429 => "0000000000000000", 13430 => "0000000000000000", 13431 => "0000000000000000", 13432 => "0000000000000000", 13433 => "0000000000000000", 13434 => "0000000000000000", 13435 => "0000000000000000", 13436 => "0000000000000000", 13437 => "0000000000000000", 13438 => "0000000000000000", 13439 => "0000000000000000", 13440 => "0000000000000000", 13441 => "0000000000000000", 13442 => "0000000000000000", 13443 => "0000000000000000", 13444 => "0000000000000000", 13445 => "0000000000000000", 13446 => "0000000000000000", 13447 => "0000000000000000", 13448 => "0000000000000000", 13449 => "0000000000000000", 13450 => "0000000000000000", 13451 => "0000000000000000", 13452 => "0000000000000000", 13453 => "0000000000000000", 13454 => "0000000000000000", 13455 => "0000000000000000", 13456 => "0000000000000000", 13457 => "0000000000000000", 13458 => "0000000000000000", 13459 => "0000000000000000", 13460 => "0000000000000000", 13461 => "0000000000000000", 13462 => "0000000000000000", 13463 => "0000000000000000", 13464 => "0000000000000000", 13465 => "0000000000000000", 13466 => "0000000000000000", 13467 => "0000000000000000", 13468 => "0000000000000000", 13469 => "0000000000000000", 13470 => "0000000000000000", 13471 => "0000000000000000", 13472 => "0000000000000000", 13473 => "0000000000000000", 13474 => "0000000000000000", 13475 => "0000000000000000", 13476 => "0000000000000000", 13477 => "0000000000000000", 13478 => "0000000000000000", 13479 => "0000000000000000", 13480 => "0000000000000000", 13481 => "0000000000000000", 13482 => "0000000000000000", 13483 => "0000000000000000", 13484 => "0000000000000000", 13485 => "0000000000000000", 13486 => "0000000000000000", 13487 => "0000000000000000", 13488 => "0000000000000000", 13489 => "0000000000000000", 13490 => "0000000000000000", 13491 => "0000000000000000", 13492 => "0000000000000000", 13493 => "0000000000000000", 13494 => "0000000000000000", 13495 => "0000000000000000", 13496 => "0000000000000000", 13497 => "0000000000000000", 13498 => "0000000000000000", 13499 => "0000000000000000", 13500 => "0000000000000000", 13501 => "0000000000000000", 13502 => "0000000000000000", 13503 => "0000000000000000", 13504 => "0000000000000000", 13505 => "0000000000000000", 13506 => "0000000000000000", 13507 => "0000000000000000", 13508 => "0000000000000000", 13509 => "0000000000000000", 13510 => "0000000000000000", 13511 => "0000000000000000", 13512 => "0000000000000000", 13513 => "0000000000000000", 13514 => "0000000000000000", 13515 => "0000000000000000", 13516 => "0000000000000000", 13517 => "0000000000000000", 13518 => "0000000000000000", 13519 => "0000000000000000", 13520 => "0000000000000000", 13521 => "0000000000000000", 13522 => "0000000000000000", 13523 => "0000000000000000", 13524 => "0000000000000000", 13525 => "0000000000000000", 13526 => "0000000000000000", 13527 => "0000000000000000", 13528 => "0000000000000000", 13529 => "0000000000000000", 13530 => "0000000000000000", 13531 => "0000000000000000", 13532 => "0000000000000000", 13533 => "0000000000000000", 13534 => "0000000000000000", 13535 => "0000000000000000", 13536 => "0000000000000000", 13537 => "0000000000000000", 13538 => "0000000000000000", 13539 => "0000000000000000", 13540 => "0000000000000000", 13541 => "0000000000000000", 13542 => "0000000000000000", 13543 => "0000000000000000", 13544 => "0000000000000000", 13545 => "0000000000000000", 13546 => "0000000000000000", 13547 => "0000000000000000", 13548 => "0000000000000000", 13549 => "0000000000000000", 13550 => "0000000000000000", 13551 => "0000000000000000", 13552 => "0000000000000000", 13553 => "0000000000000000", 13554 => "0000000000000000", 13555 => "0000000000000000", 13556 => "0000000000000000", 13557 => "0000000000000000", 13558 => "0000000000000000", 13559 => "0000000000000000", 13560 => "0000000000000000", 13561 => "0000000000000000", 13562 => "0000000000000000", 13563 => "0000000000000000", 13564 => "0000000000000000", 13565 => "0000000000000000", 13566 => "0000000000000000", 13567 => "0000000000000000", 13568 => "0000000000000000", 13569 => "0000000000000000", 13570 => "0000000000000000", 13571 => "0000000000000000", 13572 => "0000000000000000", 13573 => "0000000000000000", 13574 => "0000000000000000", 13575 => "0000000000000000", 13576 => "0000000000000000", 13577 => "0000000000000000", 13578 => "0000000000000000", 13579 => "0000000000000000", 13580 => "0000000000000000", 13581 => "0000000000000000", 13582 => "0000000000000000", 13583 => "0000000000000000", 13584 => "0000000000000000", 13585 => "0000000000000000", 13586 => "0000000000000000", 13587 => "0000000000000000", 13588 => "0000000000000000", 13589 => "0000000000000000", 13590 => "0000000000000000", 13591 => "0000000000000000", 13592 => "0000000000000000", 13593 => "0000000000000000", 13594 => "0000000000000000", 13595 => "0000000000000000", 13596 => "0000000000000000", 13597 => "0000000000000000", 13598 => "0000000000000000", 13599 => "0000000000000000", 13600 => "0000000000000000", 13601 => "0000000000000000", 13602 => "0000000000000000", 13603 => "0000000000000000", 13604 => "0000000000000000", 13605 => "0000000000000000", 13606 => "0000000000000000", 13607 => "0000000000000000", 13608 => "0000000000000000", 13609 => "0000000000000000", 13610 => "0000000000000000", 13611 => "0000000000000000", 13612 => "0000000000000000", 13613 => "0000000000000000", 13614 => "0000000000000000", 13615 => "0000000000000000", 13616 => "0000000000000000", 13617 => "0000000000000000", 13618 => "0000000000000000", 13619 => "0000000000000000", 13620 => "0000000000000000", 13621 => "0000000000000000", 13622 => "0000000000000000", 13623 => "0000000000000000", 13624 => "0000000000000000", 13625 => "0000000000000000", 13626 => "0000000000000000", 13627 => "0000000000000000", 13628 => "0000000000000000", 13629 => "0000000000000000", 13630 => "0000000000000000", 13631 => "0000000000000000", 13632 => "0000000000000000", 13633 => "0000000000000000", 13634 => "0000000000000000", 13635 => "0000000000000000", 13636 => "0000000000000000", 13637 => "0000000000000000", 13638 => "0000000000000000", 13639 => "0000000000000000", 13640 => "0000000000000000", 13641 => "0000000000000000", 13642 => "0000000000000000", 13643 => "0000000000000000", 13644 => "0000000000000000", 13645 => "0000000000000000", 13646 => "0000000000000000", 13647 => "0000000000000000", 13648 => "0000000000000000", 13649 => "0000000000000000", 13650 => "0000000000000000", 13651 => "0000000000000000", 13652 => "0000000000000000", 13653 => "0000000000000000", 13654 => "0000000000000000", 13655 => "0000000000000000", 13656 => "0000000000000000", 13657 => "0000000000000000", 13658 => "0000000000000000", 13659 => "0000000000000000", 13660 => "0000000000000000", 13661 => "0000000000000000", 13662 => "0000000000000000", 13663 => "0000000000000000", 13664 => "0000000000000000", 13665 => "0000000000000000", 13666 => "0000000000000000", 13667 => "0000000000000000", 13668 => "0000000000000000", 13669 => "0000000000000000", 13670 => "0000000000000000", 13671 => "0000000000000000", 13672 => "0000000000000000", 13673 => "0000000000000000", 13674 => "0000000000000000", 13675 => "0000000000000000", 13676 => "0000000000000000", 13677 => "0000000000000000", 13678 => "0000000000000000", 13679 => "0000000000000000", 13680 => "0000000000000000", 13681 => "0000000000000000", 13682 => "0000000000000000", 13683 => "0000000000000000", 13684 => "0000000000000000", 13685 => "0000000000000000", 13686 => "0000000000000000", 13687 => "0000000000000000", 13688 => "0000000000000000", 13689 => "0000000000000000", 13690 => "0000000000000000", 13691 => "0000000000000000", 13692 => "0000000000000000", 13693 => "0000000000000000", 13694 => "0000000000000000", 13695 => "0000000000000000", 13696 => "0000000000000000", 13697 => "0000000000000000", 13698 => "0000000000000000", 13699 => "0000000000000000", 13700 => "0000000000000000", 13701 => "0000000000000000", 13702 => "0000000000000000", 13703 => "0000000000000000", 13704 => "0000000000000000", 13705 => "0000000000000000", 13706 => "0000000000000000", 13707 => "0000000000000000", 13708 => "0000000000000000", 13709 => "0000000000000000", 13710 => "0000000000000000", 13711 => "0000000000000000", 13712 => "0000000000000000", 13713 => "0000000000000000", 13714 => "0000000000000000", 13715 => "0000000000000000", 13716 => "0000000000000000", 13717 => "0000000000000000", 13718 => "0000000000000000", 13719 => "0000000000000000", 13720 => "0000000000000000", 13721 => "0000000000000000", 13722 => "0000000000000000", 13723 => "0000000000000000", 13724 => "0000000000000000", 13725 => "0000000000000000", 13726 => "0000000000000000", 13727 => "0000000000000000", 13728 => "0000000000000000", 13729 => "0000000000000000", 13730 => "0000000000000000", 13731 => "0000000000000000", 13732 => "0000000000000000", 13733 => "0000000000000000", 13734 => "0000000000000000", 13735 => "0000000000000000", 13736 => "0000000000000000", 13737 => "0000000000000000", 13738 => "0000000000000000", 13739 => "0000000000000000", 13740 => "0000000000000000", 13741 => "0000000000000000", 13742 => "0000000000000000", 13743 => "0000000000000000", 13744 => "0000000000000000", 13745 => "0000000000000000", 13746 => "0000000000000000", 13747 => "0000000000000000", 13748 => "0000000000000000", 13749 => "0000000000000000", 13750 => "0000000000000000", 13751 => "0000000000000000", 13752 => "0000000000000000", 13753 => "0000000000000000", 13754 => "0000000000000000", 13755 => "0000000000000000", 13756 => "0000000000000000", 13757 => "0000000000000000", 13758 => "0000000000000000", 13759 => "0000000000000000", 13760 => "0000000000000000", 13761 => "0000000000000000", 13762 => "0000000000000000", 13763 => "0000000000000000", 13764 => "0000000000000000", 13765 => "0000000000000000", 13766 => "0000000000000000", 13767 => "0000000000000000", 13768 => "0000000000000000", 13769 => "0000000000000000", 13770 => "0000000000000000", 13771 => "0000000000000000", 13772 => "0000000000000000", 13773 => "0000000000000000", 13774 => "0000000000000000", 13775 => "0000000000000000", 13776 => "0000000000000000", 13777 => "0000000000000000", 13778 => "0000000000000000", 13779 => "0000000000000000", 13780 => "0000000000000000", 13781 => "0000000000000000", 13782 => "0000000000000000", 13783 => "0000000000000000", 13784 => "0000000000000000", 13785 => "0000000000000000", 13786 => "0000000000000000", 13787 => "0000000000000000", 13788 => "0000000000000000", 13789 => "0000000000000000", 13790 => "0000000000000000", 13791 => "0000000000000000", 13792 => "0000000000000000", 13793 => "0000000000000000", 13794 => "0000000000000000", 13795 => "0000000000000000", 13796 => "0000000000000000", 13797 => "0000000000000000", 13798 => "0000000000000000", 13799 => "0000000000000000", 13800 => "0000000000000000", 13801 => "0000000000000000", 13802 => "0000000000000000", 13803 => "0000000000000000", 13804 => "0000000000000000", 13805 => "0000000000000000", 13806 => "0000000000000000", 13807 => "0000000000000000", 13808 => "0000000000000000", 13809 => "0000000000000000", 13810 => "0000000000000000", 13811 => "0000000000000000", 13812 => "0000000000000000", 13813 => "0000000000000000", 13814 => "0000000000000000", 13815 => "0000000000000000", 13816 => "0000000000000000", 13817 => "0000000000000000", 13818 => "0000000000000000", 13819 => "0000000000000000", 13820 => "0000000000000000", 13821 => "0000000000000000", 13822 => "0000000000000000", 13823 => "0000000000000000", 13824 => "0000000000000000", 13825 => "0000000000000000", 13826 => "0000000000000000", 13827 => "0000000000000000", 13828 => "0000000000000000", 13829 => "0000000000000000", 13830 => "0000000000000000", 13831 => "0000000000000000", 13832 => "0000000000000000", 13833 => "0000000000000000", 13834 => "0000000000000000", 13835 => "0000000000000000", 13836 => "0000000000000000", 13837 => "0000000000000000", 13838 => "0000000000000000", 13839 => "0000000000000000", 13840 => "0000000000000000", 13841 => "0000000000000000", 13842 => "0000000000000000", 13843 => "0000000000000000", 13844 => "0000000000000000", 13845 => "0000000000000000", 13846 => "0000000000000000", 13847 => "0000000000000000", 13848 => "0000000000000000", 13849 => "0000000000000000", 13850 => "0000000000000000", 13851 => "0000000000000000", 13852 => "0000000000000000", 13853 => "0000000000000000", 13854 => "0000000000000000", 13855 => "0000000000000000", 13856 => "0000000000000000", 13857 => "0000000000000000", 13858 => "0000000000000000", 13859 => "0000000000000000", 13860 => "0000000000000000", 13861 => "0000000000000000", 13862 => "0000000000000000", 13863 => "0000000000000000", 13864 => "0000000000000000", 13865 => "0000000000000000", 13866 => "0000000000000000", 13867 => "0000000000000000", 13868 => "0000000000000000", 13869 => "0000000000000000", 13870 => "0000000000000000", 13871 => "0000000000000000", 13872 => "0000000000000000", 13873 => "0000000000000000", 13874 => "0000000000000000", 13875 => "0000000000000000", 13876 => "0000000000000000", 13877 => "0000000000000000", 13878 => "0000000000000000", 13879 => "0000000000000000", 13880 => "0000000000000000", 13881 => "0000000000000000", 13882 => "0000000000000000", 13883 => "0000000000000000", 13884 => "0000000000000000", 13885 => "0000000000000000", 13886 => "0000000000000000", 13887 => "0000000000000000", 13888 => "0000000000000000", 13889 => "0000000000000000", 13890 => "0000000000000000", 13891 => "0000000000000000", 13892 => "0000000000000000", 13893 => "0000000000000000", 13894 => "0000000000000000", 13895 => "0000000000000000", 13896 => "0000000000000000", 13897 => "0000000000000000", 13898 => "0000000000000000", 13899 => "0000000000000000", 13900 => "0000000000000000", 13901 => "0000000000000000", 13902 => "0000000000000000", 13903 => "0000000000000000", 13904 => "0000000000000000", 13905 => "0000000000000000", 13906 => "0000000000000000", 13907 => "0000000000000000", 13908 => "0000000000000000", 13909 => "0000000000000000", 13910 => "0000000000000000", 13911 => "0000000000000000", 13912 => "0000000000000000", 13913 => "0000000000000000", 13914 => "0000000000000000", 13915 => "0000000000000000", 13916 => "0000000000000000", 13917 => "0000000000000000", 13918 => "0000000000000000", 13919 => "0000000000000000", 13920 => "0000000000000000", 13921 => "0000000000000000", 13922 => "0000000000000000", 13923 => "0000000000000000", 13924 => "0000000000000000", 13925 => "0000000000000000", 13926 => "0000000000000000", 13927 => "0000000000000000", 13928 => "0000000000000000", 13929 => "0000000000000000", 13930 => "0000000000000000", 13931 => "0000000000000000", 13932 => "0000000000000000", 13933 => "0000000000000000", 13934 => "0000000000000000", 13935 => "0000000000000000", 13936 => "0000000000000000", 13937 => "0000000000000000", 13938 => "0000000000000000", 13939 => "0000000000000000", 13940 => "0000000000000000", 13941 => "0000000000000000", 13942 => "0000000000000000", 13943 => "0000000000000000", 13944 => "0000000000000000", 13945 => "0000000000000000", 13946 => "0000000000000000", 13947 => "0000000000000000", 13948 => "0000000000000000", 13949 => "0000000000000000", 13950 => "0000000000000000", 13951 => "0000000000000000", 13952 => "0000000000000000", 13953 => "0000000000000000", 13954 => "0000000000000000", 13955 => "0000000000000000", 13956 => "0000000000000000", 13957 => "0000000000000000", 13958 => "0000000000000000", 13959 => "0000000000000000", 13960 => "0000000000000000", 13961 => "0000000000000000", 13962 => "0000000000000000", 13963 => "0000000000000000", 13964 => "0000000000000000", 13965 => "0000000000000000", 13966 => "0000000000000000", 13967 => "0000000000000000", 13968 => "0000000000000000", 13969 => "0000000000000000", 13970 => "0000000000000000", 13971 => "0000000000000000", 13972 => "0000000000000000", 13973 => "0000000000000000", 13974 => "0000000000000000", 13975 => "0000000000000000", 13976 => "0000000000000000", 13977 => "0000000000000000", 13978 => "0000000000000000", 13979 => "0000000000000000", 13980 => "0000000000000000", 13981 => "0000000000000000", 13982 => "0000000000000000", 13983 => "0000000000000000", 13984 => "0000000000000000", 13985 => "0000000000000000", 13986 => "0000000000000000", 13987 => "0000000000000000", 13988 => "0000000000000000", 13989 => "0000000000000000", 13990 => "0000000000000000", 13991 => "0000000000000000", 13992 => "0000000000000000", 13993 => "0000000000000000", 13994 => "0000000000000000", 13995 => "0000000000000000", 13996 => "0000000000000000", 13997 => "0000000000000000", 13998 => "0000000000000000", 13999 => "0000000000000000", 14000 => "0000000000000000", 14001 => "0000000000000000", 14002 => "0000000000000000", 14003 => "0000000000000000", 14004 => "0000000000000000", 14005 => "0000000000000000", 14006 => "0000000000000000", 14007 => "0000000000000000", 14008 => "0000000000000000", 14009 => "0000000000000000", 14010 => "0000000000000000", 14011 => "0000000000000000", 14012 => "0000000000000000", 14013 => "0000000000000000", 14014 => "0000000000000000", 14015 => "0000000000000000", 14016 => "0000000000000000", 14017 => "0000000000000000", 14018 => "0000000000000000", 14019 => "0000000000000000", 14020 => "0000000000000000", 14021 => "0000000000000000", 14022 => "0000000000000000", 14023 => "0000000000000000", 14024 => "0000000000000000", 14025 => "0000000000000000", 14026 => "0000000000000000", 14027 => "0000000000000000", 14028 => "0000000000000000", 14029 => "0000000000000000", 14030 => "0000000000000000", 14031 => "0000000000000000", 14032 => "0000000000000000", 14033 => "0000000000000000", 14034 => "0000000000000000", 14035 => "0000000000000000", 14036 => "0000000000000000", 14037 => "0000000000000000", 14038 => "0000000000000000", 14039 => "0000000000000000", 14040 => "0000000000000000", 14041 => "0000000000000000", 14042 => "0000000000000000", 14043 => "0000000000000000", 14044 => "0000000000000000", 14045 => "0000000000000000", 14046 => "0000000000000000", 14047 => "0000000000000000", 14048 => "0000000000000000", 14049 => "0000000000000000", 14050 => "0000000000000000", 14051 => "0000000000000000", 14052 => "0000000000000000", 14053 => "0000000000000000", 14054 => "0000000000000000", 14055 => "0000000000000000", 14056 => "0000000000000000", 14057 => "0000000000000000", 14058 => "0000000000000000", 14059 => "0000000000000000", 14060 => "0000000000000000", 14061 => "0000000000000000", 14062 => "0000000000000000", 14063 => "0000000000000000", 14064 => "0000000000000000", 14065 => "0000000000000000", 14066 => "0000000000000000", 14067 => "0000000000000000", 14068 => "0000000000000000", 14069 => "0000000000000000", 14070 => "0000000000000000", 14071 => "0000000000000000", 14072 => "0000000000000000", 14073 => "0000000000000000", 14074 => "0000000000000000", 14075 => "0000000000000000", 14076 => "0000000000000000", 14077 => "0000000000000000", 14078 => "0000000000000000", 14079 => "0000000000000000", 14080 => "0000000000000000", 14081 => "0000000000000000", 14082 => "0000000000000000", 14083 => "0000000000000000", 14084 => "0000000000000000", 14085 => "0000000000000000", 14086 => "0000000000000000", 14087 => "0000000000000000", 14088 => "0000000000000000", 14089 => "0000000000000000", 14090 => "0000000000000000", 14091 => "0000000000000000", 14092 => "0000000000000000", 14093 => "0000000000000000", 14094 => "0000000000000000", 14095 => "0000000000000000", 14096 => "0000000000000000", 14097 => "0000000000000000", 14098 => "0000000000000000", 14099 => "0000000000000000", 14100 => "0000000000000000", 14101 => "0000000000000000", 14102 => "0000000000000000", 14103 => "0000000000000000", 14104 => "0000000000000000", 14105 => "0000000000000000", 14106 => "0000000000000000", 14107 => "0000000000000000", 14108 => "0000000000000000", 14109 => "0000000000000000", 14110 => "0000000000000000", 14111 => "0000000000000000", 14112 => "0000000000000000", 14113 => "0000000000000000", 14114 => "0000000000000000", 14115 => "0000000000000000", 14116 => "0000000000000000", 14117 => "0000000000000000", 14118 => "0000000000000000", 14119 => "0000000000000000", 14120 => "0000000000000000", 14121 => "0000000000000000", 14122 => "0000000000000000", 14123 => "0000000000000000", 14124 => "0000000000000000", 14125 => "0000000000000000", 14126 => "0000000000000000", 14127 => "0000000000000000", 14128 => "0000000000000000", 14129 => "0000000000000000", 14130 => "0000000000000000", 14131 => "0000000000000000", 14132 => "0000000000000000", 14133 => "0000000000000000", 14134 => "0000000000000000", 14135 => "0000000000000000", 14136 => "0000000000000000", 14137 => "0000000000000000", 14138 => "0000000000000000", 14139 => "0000000000000000", 14140 => "0000000000000000", 14141 => "0000000000000000", 14142 => "0000000000000000", 14143 => "0000000000000000", 14144 => "0000000000000000", 14145 => "0000000000000000", 14146 => "0000000000000000", 14147 => "0000000000000000", 14148 => "0000000000000000", 14149 => "0000000000000000", 14150 => "0000000000000000", 14151 => "0000000000000000", 14152 => "0000000000000000", 14153 => "0000000000000000", 14154 => "0000000000000000", 14155 => "0000000000000000", 14156 => "0000000000000000", 14157 => "0000000000000000", 14158 => "0000000000000000", 14159 => "0000000000000000", 14160 => "0000000000000000", 14161 => "0000000000000000", 14162 => "0000000000000000", 14163 => "0000000000000000", 14164 => "0000000000000000", 14165 => "0000000000000000", 14166 => "0000000000000000", 14167 => "0000000000000000", 14168 => "0000000000000000", 14169 => "0000000000000000", 14170 => "0000000000000000", 14171 => "0000000000000000", 14172 => "0000000000000000", 14173 => "0000000000000000", 14174 => "0000000000000000", 14175 => "0000000000000000", 14176 => "0000000000000000", 14177 => "0000000000000000", 14178 => "0000000000000000", 14179 => "0000000000000000", 14180 => "0000000000000000", 14181 => "0000000000000000", 14182 => "0000000000000000", 14183 => "0000000000000000", 14184 => "0000000000000000", 14185 => "0000000000000000", 14186 => "0000000000000000", 14187 => "0000000000000000", 14188 => "0000000000000000", 14189 => "0000000000000000", 14190 => "0000000000000000", 14191 => "0000000000000000", 14192 => "0000000000000000", 14193 => "0000000000000000", 14194 => "0000000000000000", 14195 => "0000000000000000", 14196 => "0000000000000000", 14197 => "0000000000000000", 14198 => "0000000000000000", 14199 => "0000000000000000", 14200 => "0000000000000000", 14201 => "0000000000000000", 14202 => "0000000000000000", 14203 => "0000000000000000", 14204 => "0000000000000000", 14205 => "0000000000000000", 14206 => "0000000000000000", 14207 => "0000000000000000", 14208 => "0000000000000000", 14209 => "0000000000000000", 14210 => "0000000000000000", 14211 => "0000000000000000", 14212 => "0000000000000000", 14213 => "0000000000000000", 14214 => "0000000000000000", 14215 => "0000000000000000", 14216 => "0000000000000000", 14217 => "0000000000000000", 14218 => "0000000000000000", 14219 => "0000000000000000", 14220 => "0000000000000000", 14221 => "0000000000000000", 14222 => "0000000000000000", 14223 => "0000000000000000", 14224 => "0000000000000000", 14225 => "0000000000000000", 14226 => "0000000000000000", 14227 => "0000000000000000", 14228 => "0000000000000000", 14229 => "0000000000000000", 14230 => "0000000000000000", 14231 => "0000000000000000", 14232 => "0000000000000000", 14233 => "0000000000000000", 14234 => "0000000000000000", 14235 => "0000000000000000", 14236 => "0000000000000000", 14237 => "0000000000000000", 14238 => "0000000000000000", 14239 => "0000000000000000", 14240 => "0000000000000000", 14241 => "0000000000000000", 14242 => "0000000000000000", 14243 => "0000000000000000", 14244 => "0000000000000000", 14245 => "0000000000000000", 14246 => "0000000000000000", 14247 => "0000000000000000", 14248 => "0000000000000000", 14249 => "0000000000000000", 14250 => "0000000000000000", 14251 => "0000000000000000", 14252 => "0000000000000000", 14253 => "0000000000000000", 14254 => "0000000000000000", 14255 => "0000000000000000", 14256 => "0000000000000000", 14257 => "0000000000000000", 14258 => "0000000000000000", 14259 => "0000000000000000", 14260 => "0000000000000000", 14261 => "0000000000000000", 14262 => "0000000000000000", 14263 => "0000000000000000", 14264 => "0000000000000000", 14265 => "0000000000000000", 14266 => "0000000000000000", 14267 => "0000000000000000", 14268 => "0000000000000000", 14269 => "0000000000000000", 14270 => "0000000000000000", 14271 => "0000000000000000", 14272 => "0000000000000000", 14273 => "0000000000000000", 14274 => "0000000000000000", 14275 => "0000000000000000", 14276 => "0000000000000000", 14277 => "0000000000000000", 14278 => "0000000000000000", 14279 => "0000000000000000", 14280 => "0000000000000000", 14281 => "0000000000000000", 14282 => "0000000000000000", 14283 => "0000000000000000", 14284 => "0000000000000000", 14285 => "0000000000000000", 14286 => "0000000000000000", 14287 => "0000000000000000", 14288 => "0000000000000000", 14289 => "0000000000000000", 14290 => "0000000000000000", 14291 => "0000000000000000", 14292 => "0000000000000000", 14293 => "0000000000000000", 14294 => "0000000000000000", 14295 => "0000000000000000", 14296 => "0000000000000000", 14297 => "0000000000000000", 14298 => "0000000000000000", 14299 => "0000000000000000", 14300 => "0000000000000000", 14301 => "0000000000000000", 14302 => "0000000000000000", 14303 => "0000000000000000", 14304 => "0000000000000000", 14305 => "0000000000000000", 14306 => "0000000000000000", 14307 => "0000000000000000", 14308 => "0000000000000000", 14309 => "0000000000000000", 14310 => "0000000000000000", 14311 => "0000000000000000", 14312 => "0000000000000000", 14313 => "0000000000000000", 14314 => "0000000000000000", 14315 => "0000000000000000", 14316 => "0000000000000000", 14317 => "0000000000000000", 14318 => "0000000000000000", 14319 => "0000000000000000", 14320 => "0000000000000000", 14321 => "0000000000000000", 14322 => "0000000000000000", 14323 => "0000000000000000", 14324 => "0000000000000000", 14325 => "0000000000000000", 14326 => "0000000000000000", 14327 => "0000000000000000", 14328 => "0000000000000000", 14329 => "0000000000000000", 14330 => "0000000000000000", 14331 => "0000000000000000", 14332 => "0000000000000000", 14333 => "0000000000000000", 14334 => "0000000000000000", 14335 => "0000000000000000", 14336 => "0000000000000000", 14337 => "0000000000000000", 14338 => "0000000000000000", 14339 => "0000000000000000", 14340 => "0000000000000000", 14341 => "0000000000000000", 14342 => "0000000000000000", 14343 => "0000000000000000", 14344 => "0000000000000000", 14345 => "0000000000000000", 14346 => "0000000000000000", 14347 => "0000000000000000", 14348 => "0000000000000000", 14349 => "0000000000000000", 14350 => "0000000000000000", 14351 => "0000000000000000", 14352 => "0000000000000000", 14353 => "0000000000000000", 14354 => "0000000000000000", 14355 => "0000000000000000", 14356 => "0000000000000000", 14357 => "0000000000000000", 14358 => "0000000000000000", 14359 => "0000000000000000", 14360 => "0000000000000000", 14361 => "0000000000000000", 14362 => "0000000000000000", 14363 => "0000000000000000", 14364 => "0000000000000000", 14365 => "0000000000000000", 14366 => "0000000000000000", 14367 => "0000000000000000", 14368 => "0000000000000000", 14369 => "0000000000000000", 14370 => "0000000000000000", 14371 => "0000000000000000", 14372 => "0000000000000000", 14373 => "0000000000000000", 14374 => "0000000000000000", 14375 => "0000000000000000", 14376 => "0000000000000000", 14377 => "0000000000000000", 14378 => "0000000000000000", 14379 => "0000000000000000", 14380 => "0000000000000000", 14381 => "0000000000000000", 14382 => "0000000000000000", 14383 => "0000000000000000", 14384 => "0000000000000000", 14385 => "0000000000000000", 14386 => "0000000000000000", 14387 => "0000000000000000", 14388 => "0000000000000000", 14389 => "0000000000000000", 14390 => "0000000000000000", 14391 => "0000000000000000", 14392 => "0000000000000000", 14393 => "0000000000000000", 14394 => "0000000000000000", 14395 => "0000000000000000", 14396 => "0000000000000000", 14397 => "0000000000000000", 14398 => "0000000000000000", 14399 => "0000000000000000", 14400 => "0000000000000000", 14401 => "0000000000000000", 14402 => "0000000000000000", 14403 => "0000000000000000", 14404 => "0000000000000000", 14405 => "0000000000000000", 14406 => "0000000000000000", 14407 => "0000000000000000", 14408 => "0000000000000000", 14409 => "0000000000000000", 14410 => "0000000000000000", 14411 => "0000000000000000", 14412 => "0000000000000000", 14413 => "0000000000000000", 14414 => "0000000000000000", 14415 => "0000000000000000", 14416 => "0000000000000000", 14417 => "0000000000000000", 14418 => "0000000000000000", 14419 => "0000000000000000", 14420 => "0000000000000000", 14421 => "0000000000000000", 14422 => "0000000000000000", 14423 => "0000000000000000", 14424 => "0000000000000000", 14425 => "0000000000000000", 14426 => "0000000000000000", 14427 => "0000000000000000", 14428 => "0000000000000000", 14429 => "0000000000000000", 14430 => "0000000000000000", 14431 => "0000000000000000", 14432 => "0000000000000000", 14433 => "0000000000000000", 14434 => "0000000000000000", 14435 => "0000000000000000", 14436 => "0000000000000000", 14437 => "0000000000000000", 14438 => "0000000000000000", 14439 => "0000000000000000", 14440 => "0000000000000000", 14441 => "0000000000000000", 14442 => "0000000000000000", 14443 => "0000000000000000", 14444 => "0000000000000000", 14445 => "0000000000000000", 14446 => "0000000000000000", 14447 => "0000000000000000", 14448 => "0000000000000000", 14449 => "0000000000000000", 14450 => "0000000000000000", 14451 => "0000000000000000", 14452 => "0000000000000000", 14453 => "0000000000000000", 14454 => "0000000000000000", 14455 => "0000000000000000", 14456 => "0000000000000000", 14457 => "0000000000000000", 14458 => "0000000000000000", 14459 => "0000000000000000", 14460 => "0000000000000000", 14461 => "0000000000000000", 14462 => "0000000000000000", 14463 => "0000000000000000", 14464 => "0000000000000000", 14465 => "0000000000000000", 14466 => "0000000000000000", 14467 => "0000000000000000", 14468 => "0000000000000000", 14469 => "0000000000000000", 14470 => "0000000000000000", 14471 => "0000000000000000", 14472 => "0000000000000000", 14473 => "0000000000000000", 14474 => "0000000000000000", 14475 => "0000000000000000", 14476 => "0000000000000000", 14477 => "0000000000000000", 14478 => "0000000000000000", 14479 => "0000000000000000", 14480 => "0000000000000000", 14481 => "0000000000000000", 14482 => "0000000000000000", 14483 => "0000000000000000", 14484 => "0000000000000000", 14485 => "0000000000000000", 14486 => "0000000000000000", 14487 => "0000000000000000", 14488 => "0000000000000000", 14489 => "0000000000000000", 14490 => "0000000000000000", 14491 => "0000000000000000", 14492 => "0000000000000000", 14493 => "0000000000000000", 14494 => "0000000000000000", 14495 => "0000000000000000", 14496 => "0000000000000000", 14497 => "0000000000000000", 14498 => "0000000000000000", 14499 => "0000000000000000", 14500 => "0000000000000000", 14501 => "0000000000000000", 14502 => "0000000000000000", 14503 => "0000000000000000", 14504 => "0000000000000000", 14505 => "0000000000000000", 14506 => "0000000000000000", 14507 => "0000000000000000", 14508 => "0000000000000000", 14509 => "0000000000000000", 14510 => "0000000000000000", 14511 => "0000000000000000", 14512 => "0000000000000000", 14513 => "0000000000000000", 14514 => "0000000000000000", 14515 => "0000000000000000", 14516 => "0000000000000000", 14517 => "0000000000000000", 14518 => "0000000000000000", 14519 => "0000000000000000", 14520 => "0000000000000000", 14521 => "0000000000000000", 14522 => "0000000000000000", 14523 => "0000000000000000", 14524 => "0000000000000000", 14525 => "0000000000000000", 14526 => "0000000000000000", 14527 => "0000000000000000", 14528 => "0000000000000000", 14529 => "0000000000000000", 14530 => "0000000000000000", 14531 => "0000000000000000", 14532 => "0000000000000000", 14533 => "0000000000000000", 14534 => "0000000000000000", 14535 => "0000000000000000", 14536 => "0000000000000000", 14537 => "0000000000000000", 14538 => "0000000000000000", 14539 => "0000000000000000", 14540 => "0000000000000000", 14541 => "0000000000000000", 14542 => "0000000000000000", 14543 => "0000000000000000", 14544 => "0000000000000000", 14545 => "0000000000000000", 14546 => "0000000000000000", 14547 => "0000000000000000", 14548 => "0000000000000000", 14549 => "0000000000000000", 14550 => "0000000000000000", 14551 => "0000000000000000", 14552 => "0000000000000000", 14553 => "0000000000000000", 14554 => "0000000000000000", 14555 => "0000000000000000", 14556 => "0000000000000000", 14557 => "0000000000000000", 14558 => "0000000000000000", 14559 => "0000000000000000", 14560 => "0000000000000000", 14561 => "0000000000000000", 14562 => "0000000000000000", 14563 => "0000000000000000", 14564 => "0000000000000000", 14565 => "0000000000000000", 14566 => "0000000000000000", 14567 => "0000000000000000", 14568 => "0000000000000000", 14569 => "0000000000000000", 14570 => "0000000000000000", 14571 => "0000000000000000", 14572 => "0000000000000000", 14573 => "0000000000000000", 14574 => "0000000000000000", 14575 => "0000000000000000", 14576 => "0000000000000000", 14577 => "0000000000000000", 14578 => "0000000000000000", 14579 => "0000000000000000", 14580 => "0000000000000000", 14581 => "0000000000000000", 14582 => "0000000000000000", 14583 => "0000000000000000", 14584 => "0000000000000000", 14585 => "0000000000000000", 14586 => "0000000000000000", 14587 => "0000000000000000", 14588 => "0000000000000000", 14589 => "0000000000000000", 14590 => "0000000000000000", 14591 => "0000000000000000", 14592 => "0000000000000000", 14593 => "0000000000000000", 14594 => "0000000000000000", 14595 => "0000000000000000", 14596 => "0000000000000000", 14597 => "0000000000000000", 14598 => "0000000000000000", 14599 => "0000000000000000", 14600 => "0000000000000000", 14601 => "0000000000000000", 14602 => "0000000000000000", 14603 => "0000000000000000", 14604 => "0000000000000000", 14605 => "0000000000000000", 14606 => "0000000000000000", 14607 => "0000000000000000", 14608 => "0000000000000000", 14609 => "0000000000000000", 14610 => "0000000000000000", 14611 => "0000000000000000", 14612 => "0000000000000000", 14613 => "0000000000000000", 14614 => "0000000000000000", 14615 => "0000000000000000", 14616 => "0000000000000000", 14617 => "0000000000000000", 14618 => "0000000000000000", 14619 => "0000000000000000", 14620 => "0000000000000000", 14621 => "0000000000000000", 14622 => "0000000000000000", 14623 => "0000000000000000", 14624 => "0000000000000000", 14625 => "0000000000000000", 14626 => "0000000000000000", 14627 => "0000000000000000", 14628 => "0000000000000000", 14629 => "0000000000000000", 14630 => "0000000000000000", 14631 => "0000000000000000", 14632 => "0000000000000000", 14633 => "0000000000000000", 14634 => "0000000000000000", 14635 => "0000000000000000", 14636 => "0000000000000000", 14637 => "0000000000000000", 14638 => "0000000000000000", 14639 => "0000000000000000", 14640 => "0000000000000000", 14641 => "0000000000000000", 14642 => "0000000000000000", 14643 => "0000000000000000", 14644 => "0000000000000000", 14645 => "0000000000000000", 14646 => "0000000000000000", 14647 => "0000000000000000", 14648 => "0000000000000000", 14649 => "0000000000000000", 14650 => "0000000000000000", 14651 => "0000000000000000", 14652 => "0000000000000000", 14653 => "0000000000000000", 14654 => "0000000000000000", 14655 => "0000000000000000", 14656 => "0000000000000000", 14657 => "0000000000000000", 14658 => "0000000000000000", 14659 => "0000000000000000", 14660 => "0000000000000000", 14661 => "0000000000000000", 14662 => "0000000000000000", 14663 => "0000000000000000", 14664 => "0000000000000000", 14665 => "0000000000000000", 14666 => "0000000000000000", 14667 => "0000000000000000", 14668 => "0000000000000000", 14669 => "0000000000000000", 14670 => "0000000000000000", 14671 => "0000000000000000", 14672 => "0000000000000000", 14673 => "0000000000000000", 14674 => "0000000000000000", 14675 => "0000000000000000", 14676 => "0000000000000000", 14677 => "0000000000000000", 14678 => "0000000000000000", 14679 => "0000000000000000", 14680 => "0000000000000000", 14681 => "0000000000000000", 14682 => "0000000000000000", 14683 => "0000000000000000", 14684 => "0000000000000000", 14685 => "0000000000000000", 14686 => "0000000000000000", 14687 => "0000000000000000", 14688 => "0000000000000000", 14689 => "0000000000000000", 14690 => "0000000000000000", 14691 => "0000000000000000", 14692 => "0000000000000000", 14693 => "0000000000000000", 14694 => "0000000000000000", 14695 => "0000000000000000", 14696 => "0000000000000000", 14697 => "0000000000000000", 14698 => "0000000000000000", 14699 => "0000000000000000", 14700 => "0000000000000000", 14701 => "0000000000000000", 14702 => "0000000000000000", 14703 => "0000000000000000", 14704 => "0000000000000000", 14705 => "0000000000000000", 14706 => "0000000000000000", 14707 => "0000000000000000", 14708 => "0000000000000000", 14709 => "0000000000000000", 14710 => "0000000000000000", 14711 => "0000000000000000", 14712 => "0000000000000000", 14713 => "0000000000000000", 14714 => "0000000000000000", 14715 => "0000000000000000", 14716 => "0000000000000000", 14717 => "0000000000000000", 14718 => "0000000000000000", 14719 => "0000000000000000", 14720 => "0000000000000000", 14721 => "0000000000000000", 14722 => "0000000000000000", 14723 => "0000000000000000", 14724 => "0000000000000000", 14725 => "0000000000000000", 14726 => "0000000000000000", 14727 => "0000000000000000", 14728 => "0000000000000000", 14729 => "0000000000000000", 14730 => "0000000000000000", 14731 => "0000000000000000", 14732 => "0000000000000000", 14733 => "0000000000000000", 14734 => "0000000000000000", 14735 => "0000000000000000", 14736 => "0000000000000000", 14737 => "0000000000000000", 14738 => "0000000000000000", 14739 => "0000000000000000", 14740 => "0000000000000000", 14741 => "0000000000000000", 14742 => "0000000000000000", 14743 => "0000000000000000", 14744 => "0000000000000000", 14745 => "0000000000000000", 14746 => "0000000000000000", 14747 => "0000000000000000", 14748 => "0000000000000000", 14749 => "0000000000000000", 14750 => "0000000000000000", 14751 => "0000000000000000", 14752 => "0000000000000000", 14753 => "0000000000000000", 14754 => "0000000000000000", 14755 => "0000000000000000", 14756 => "0000000000000000", 14757 => "0000000000000000", 14758 => "0000000000000000", 14759 => "0000000000000000", 14760 => "0000000000000000", 14761 => "0000000000000000", 14762 => "0000000000000000", 14763 => "0000000000000000", 14764 => "0000000000000000", 14765 => "0000000000000000", 14766 => "0000000000000000", 14767 => "0000000000000000", 14768 => "0000000000000000", 14769 => "0000000000000000", 14770 => "0000000000000000", 14771 => "0000000000000000", 14772 => "0000000000000000", 14773 => "0000000000000000", 14774 => "0000000000000000", 14775 => "0000000000000000", 14776 => "0000000000000000", 14777 => "0000000000000000", 14778 => "0000000000000000", 14779 => "0000000000000000", 14780 => "0000000000000000", 14781 => "0000000000000000", 14782 => "0000000000000000", 14783 => "0000000000000000", 14784 => "0000000000000000", 14785 => "0000000000000000", 14786 => "0000000000000000", 14787 => "0000000000000000", 14788 => "0000000000000000", 14789 => "0000000000000000", 14790 => "0000000000000000", 14791 => "0000000000000000", 14792 => "0000000000000000", 14793 => "0000000000000000", 14794 => "0000000000000000", 14795 => "0000000000000000", 14796 => "0000000000000000", 14797 => "0000000000000000", 14798 => "0000000000000000", 14799 => "0000000000000000", 14800 => "0000000000000000", 14801 => "0000000000000000", 14802 => "0000000000000000", 14803 => "0000000000000000", 14804 => "0000000000000000", 14805 => "0000000000000000", 14806 => "0000000000000000", 14807 => "0000000000000000", 14808 => "0000000000000000", 14809 => "0000000000000000", 14810 => "0000000000000000", 14811 => "0000000000000000", 14812 => "0000000000000000", 14813 => "0000000000000000", 14814 => "0000000000000000", 14815 => "0000000000000000", 14816 => "0000000000000000", 14817 => "0000000000000000", 14818 => "0000000000000000", 14819 => "0000000000000000", 14820 => "0000000000000000", 14821 => "0000000000000000", 14822 => "0000000000000000", 14823 => "0000000000000000", 14824 => "0000000000000000", 14825 => "0000000000000000", 14826 => "0000000000000000", 14827 => "0000000000000000", 14828 => "0000000000000000", 14829 => "0000000000000000", 14830 => "0000000000000000", 14831 => "0000000000000000", 14832 => "0000000000000000", 14833 => "0000000000000000", 14834 => "0000000000000000", 14835 => "0000000000000000", 14836 => "0000000000000000", 14837 => "0000000000000000", 14838 => "0000000000000000", 14839 => "0000000000000000", 14840 => "0000000000000000", 14841 => "0000000000000000", 14842 => "0000000000000000", 14843 => "0000000000000000", 14844 => "0000000000000000", 14845 => "0000000000000000", 14846 => "0000000000000000", 14847 => "0000000000000000", 14848 => "0000000000000000", 14849 => "0000000000000000", 14850 => "0000000000000000", 14851 => "0000000000000000", 14852 => "0000000000000000", 14853 => "0000000000000000", 14854 => "0000000000000000", 14855 => "0000000000000000", 14856 => "0000000000000000", 14857 => "0000000000000000", 14858 => "0000000000000000", 14859 => "0000000000000000", 14860 => "0000000000000000", 14861 => "0000000000000000", 14862 => "0000000000000000", 14863 => "0000000000000000", 14864 => "0000000000000000", 14865 => "0000000000000000", 14866 => "0000000000000000", 14867 => "0000000000000000", 14868 => "0000000000000000", 14869 => "0000000000000000", 14870 => "0000000000000000", 14871 => "0000000000000000", 14872 => "0000000000000000", 14873 => "0000000000000000", 14874 => "0000000000000000", 14875 => "0000000000000000", 14876 => "0000000000000000", 14877 => "0000000000000000", 14878 => "0000000000000000", 14879 => "0000000000000000", 14880 => "0000000000000000", 14881 => "0000000000000000", 14882 => "0000000000000000", 14883 => "0000000000000000", 14884 => "0000000000000000", 14885 => "0000000000000000", 14886 => "0000000000000000", 14887 => "0000000000000000", 14888 => "0000000000000000", 14889 => "0000000000000000", 14890 => "0000000000000000", 14891 => "0000000000000000", 14892 => "0000000000000000", 14893 => "0000000000000000", 14894 => "0000000000000000", 14895 => "0000000000000000", 14896 => "0000000000000000", 14897 => "0000000000000000", 14898 => "0000000000000000", 14899 => "0000000000000000", 14900 => "0000000000000000", 14901 => "0000000000000000", 14902 => "0000000000000000", 14903 => "0000000000000000", 14904 => "0000000000000000", 14905 => "0000000000000000", 14906 => "0000000000000000", 14907 => "0000000000000000", 14908 => "0000000000000000", 14909 => "0000000000000000", 14910 => "0000000000000000", 14911 => "0000000000000000", 14912 => "0000000000000000", 14913 => "0000000000000000", 14914 => "0000000000000000", 14915 => "0000000000000000", 14916 => "0000000000000000", 14917 => "0000000000000000", 14918 => "0000000000000000", 14919 => "0000000000000000", 14920 => "0000000000000000", 14921 => "0000000000000000", 14922 => "0000000000000000", 14923 => "0000000000000000", 14924 => "0000000000000000", 14925 => "0000000000000000", 14926 => "0000000000000000", 14927 => "0000000000000000", 14928 => "0000000000000000", 14929 => "0000000000000000", 14930 => "0000000000000000", 14931 => "0000000000000000", 14932 => "0000000000000000", 14933 => "0000000000000000", 14934 => "0000000000000000", 14935 => "0000000000000000", 14936 => "0000000000000000", 14937 => "0000000000000000", 14938 => "0000000000000000", 14939 => "0000000000000000", 14940 => "0000000000000000", 14941 => "0000000000000000", 14942 => "0000000000000000", 14943 => "0000000000000000", 14944 => "0000000000000000", 14945 => "0000000000000000", 14946 => "0000000000000000", 14947 => "0000000000000000", 14948 => "0000000000000000", 14949 => "0000000000000000", 14950 => "0000000000000000", 14951 => "0000000000000000", 14952 => "0000000000000000", 14953 => "0000000000000000", 14954 => "0000000000000000", 14955 => "0000000000000000", 14956 => "0000000000000000", 14957 => "0000000000000000", 14958 => "0000000000000000", 14959 => "0000000000000000", 14960 => "0000000000000000", 14961 => "0000000000000000", 14962 => "0000000000000000", 14963 => "0000000000000000", 14964 => "0000000000000000", 14965 => "0000000000000000", 14966 => "0000000000000000", 14967 => "0000000000000000", 14968 => "0000000000000000", 14969 => "0000000000000000", 14970 => "0000000000000000", 14971 => "0000000000000000", 14972 => "0000000000000000", 14973 => "0000000000000000", 14974 => "0000000000000000", 14975 => "0000000000000000", 14976 => "0000000000000000", 14977 => "0000000000000000", 14978 => "0000000000000000", 14979 => "0000000000000000", 14980 => "0000000000000000", 14981 => "0000000000000000", 14982 => "0000000000000000", 14983 => "0000000000000000", 14984 => "0000000000000000", 14985 => "0000000000000000", 14986 => "0000000000000000", 14987 => "0000000000000000", 14988 => "0000000000000000", 14989 => "0000000000000000", 14990 => "0000000000000000", 14991 => "0000000000000000", 14992 => "0000000000000000", 14993 => "0000000000000000", 14994 => "0000000000000000", 14995 => "0000000000000000", 14996 => "0000000000000000", 14997 => "0000000000000000", 14998 => "0000000000000000", 14999 => "0000000000000000", 15000 => "0000000000000000", 15001 => "0000000000000000", 15002 => "0000000000000000", 15003 => "0000000000000000", 15004 => "0000000000000000", 15005 => "0000000000000000", 15006 => "0000000000000000", 15007 => "0000000000000000", 15008 => "0000000000000000", 15009 => "0000000000000000", 15010 => "0000000000000000", 15011 => "0000000000000000", 15012 => "0000000000000000", 15013 => "0000000000000000", 15014 => "0000000000000000", 15015 => "0000000000000000", 15016 => "0000000000000000", 15017 => "0000000000000000", 15018 => "0000000000000000", 15019 => "0000000000000000", 15020 => "0000000000000000", 15021 => "0000000000000000", 15022 => "0000000000000000", 15023 => "0000000000000000", 15024 => "0000000000000000", 15025 => "0000000000000000", 15026 => "0000000000000000", 15027 => "0000000000000000", 15028 => "0000000000000000", 15029 => "0000000000000000", 15030 => "0000000000000000", 15031 => "0000000000000000", 15032 => "0000000000000000", 15033 => "0000000000000000", 15034 => "0000000000000000", 15035 => "0000000000000000", 15036 => "0000000000000000", 15037 => "0000000000000000", 15038 => "0000000000000000", 15039 => "0000000000000000", 15040 => "0000000000000000", 15041 => "0000000000000000", 15042 => "0000000000000000", 15043 => "0000000000000000", 15044 => "0000000000000000", 15045 => "0000000000000000", 15046 => "0000000000000000", 15047 => "0000000000000000", 15048 => "0000000000000000", 15049 => "0000000000000000", 15050 => "0000000000000000", 15051 => "0000000000000000", 15052 => "0000000000000000", 15053 => "0000000000000000", 15054 => "0000000000000000", 15055 => "0000000000000000", 15056 => "0000000000000000", 15057 => "0000000000000000", 15058 => "0000000000000000", 15059 => "0000000000000000", 15060 => "0000000000000000", 15061 => "0000000000000000", 15062 => "0000000000000000", 15063 => "0000000000000000", 15064 => "0000000000000000", 15065 => "0000000000000000", 15066 => "0000000000000000", 15067 => "0000000000000000", 15068 => "0000000000000000", 15069 => "0000000000000000", 15070 => "0000000000000000", 15071 => "0000000000000000", 15072 => "0000000000000000", 15073 => "0000000000000000", 15074 => "0000000000000000", 15075 => "0000000000000000", 15076 => "0000000000000000", 15077 => "0000000000000000", 15078 => "0000000000000000", 15079 => "0000000000000000", 15080 => "0000000000000000", 15081 => "0000000000000000", 15082 => "0000000000000000", 15083 => "0000000000000000", 15084 => "0000000000000000", 15085 => "0000000000000000", 15086 => "0000000000000000", 15087 => "0000000000000000", 15088 => "0000000000000000", 15089 => "0000000000000000", 15090 => "0000000000000000", 15091 => "0000000000000000", 15092 => "0000000000000000", 15093 => "0000000000000000", 15094 => "0000000000000000", 15095 => "0000000000000000", 15096 => "0000000000000000", 15097 => "0000000000000000", 15098 => "0000000000000000", 15099 => "0000000000000000", 15100 => "0000000000000000", 15101 => "0000000000000000", 15102 => "0000000000000000", 15103 => "0000000000000000", 15104 => "0000000000000000", 15105 => "0000000000000000", 15106 => "0000000000000000", 15107 => "0000000000000000", 15108 => "0000000000000000", 15109 => "0000000000000000", 15110 => "0000000000000000", 15111 => "0000000000000000", 15112 => "0000000000000000", 15113 => "0000000000000000", 15114 => "0000000000000000", 15115 => "0000000000000000", 15116 => "0000000000000000", 15117 => "0000000000000000", 15118 => "0000000000000000", 15119 => "0000000000000000", 15120 => "0000000000000000", 15121 => "0000000000000000", 15122 => "0000000000000000", 15123 => "0000000000000000", 15124 => "0000000000000000", 15125 => "0000000000000000", 15126 => "0000000000000000", 15127 => "0000000000000000", 15128 => "0000000000000000", 15129 => "0000000000000000", 15130 => "0000000000000000", 15131 => "0000000000000000", 15132 => "0000000000000000", 15133 => "0000000000000000", 15134 => "0000000000000000", 15135 => "0000000000000000", 15136 => "0000000000000000", 15137 => "0000000000000000", 15138 => "0000000000000000", 15139 => "0000000000000000", 15140 => "0000000000000000", 15141 => "0000000000000000", 15142 => "0000000000000000", 15143 => "0000000000000000", 15144 => "0000000000000000", 15145 => "0000000000000000", 15146 => "0000000000000000", 15147 => "0000000000000000", 15148 => "0000000000000000", 15149 => "0000000000000000", 15150 => "0000000000000000", 15151 => "0000000000000000", 15152 => "0000000000000000", 15153 => "0000000000000000", 15154 => "0000000000000000", 15155 => "0000000000000000", 15156 => "0000000000000000", 15157 => "0000000000000000", 15158 => "0000000000000000", 15159 => "0000000000000000", 15160 => "0000000000000000", 15161 => "0000000000000000", 15162 => "0000000000000000", 15163 => "0000000000000000", 15164 => "0000000000000000", 15165 => "0000000000000000", 15166 => "0000000000000000", 15167 => "0000000000000000", 15168 => "0000000000000000", 15169 => "0000000000000000", 15170 => "0000000000000000", 15171 => "0000000000000000", 15172 => "0000000000000000", 15173 => "0000000000000000", 15174 => "0000000000000000", 15175 => "0000000000000000", 15176 => "0000000000000000", 15177 => "0000000000000000", 15178 => "0000000000000000", 15179 => "0000000000000000", 15180 => "0000000000000000", 15181 => "0000000000000000", 15182 => "0000000000000000", 15183 => "0000000000000000", 15184 => "0000000000000000", 15185 => "0000000000000000", 15186 => "0000000000000000", 15187 => "0000000000000000", 15188 => "0000000000000000", 15189 => "0000000000000000", 15190 => "0000000000000000", 15191 => "0000000000000000", 15192 => "0000000000000000", 15193 => "0000000000000000", 15194 => "0000000000000000", 15195 => "0000000000000000", 15196 => "0000000000000000", 15197 => "0000000000000000", 15198 => "0000000000000000", 15199 => "0000000000000000", 15200 => "0000000000000000", 15201 => "0000000000000000", 15202 => "0000000000000000", 15203 => "0000000000000000", 15204 => "0000000000000000", 15205 => "0000000000000000", 15206 => "0000000000000000", 15207 => "0000000000000000", 15208 => "0000000000000000", 15209 => "0000000000000000", 15210 => "0000000000000000", 15211 => "0000000000000000", 15212 => "0000000000000000", 15213 => "0000000000000000", 15214 => "0000000000000000", 15215 => "0000000000000000", 15216 => "0000000000000000", 15217 => "0000000000000000", 15218 => "0000000000000000", 15219 => "0000000000000000", 15220 => "0000000000000000", 15221 => "0000000000000000", 15222 => "0000000000000000", 15223 => "0000000000000000", 15224 => "0000000000000000", 15225 => "0000000000000000", 15226 => "0000000000000000", 15227 => "0000000000000000", 15228 => "0000000000000000", 15229 => "0000000000000000", 15230 => "0000000000000000", 15231 => "0000000000000000", 15232 => "0000000000000000", 15233 => "0000000000000000", 15234 => "0000000000000000", 15235 => "0000000000000000", 15236 => "0000000000000000", 15237 => "0000000000000000", 15238 => "0000000000000000", 15239 => "0000000000000000", 15240 => "0000000000000000", 15241 => "0000000000000000", 15242 => "0000000000000000", 15243 => "0000000000000000", 15244 => "0000000000000000", 15245 => "0000000000000000", 15246 => "0000000000000000", 15247 => "0000000000000000", 15248 => "0000000000000000", 15249 => "0000000000000000", 15250 => "0000000000000000", 15251 => "0000000000000000", 15252 => "0000000000000000", 15253 => "0000000000000000", 15254 => "0000000000000000", 15255 => "0000000000000000", 15256 => "0000000000000000", 15257 => "0000000000000000", 15258 => "0000000000000000", 15259 => "0000000000000000", 15260 => "0000000000000000", 15261 => "0000000000000000", 15262 => "0000000000000000", 15263 => "0000000000000000", 15264 => "0000000000000000", 15265 => "0000000000000000", 15266 => "0000000000000000", 15267 => "0000000000000000", 15268 => "0000000000000000", 15269 => "0000000000000000", 15270 => "0000000000000000", 15271 => "0000000000000000", 15272 => "0000000000000000", 15273 => "0000000000000000", 15274 => "0000000000000000", 15275 => "0000000000000000", 15276 => "0000000000000000", 15277 => "0000000000000000", 15278 => "0000000000000000", 15279 => "0000000000000000", 15280 => "0000000000000000", 15281 => "0000000000000000", 15282 => "0000000000000000", 15283 => "0000000000000000", 15284 => "0000000000000000", 15285 => "0000000000000000", 15286 => "0000000000000000", 15287 => "0000000000000000", 15288 => "0000000000000000", 15289 => "0000000000000000", 15290 => "0000000000000000", 15291 => "0000000000000000", 15292 => "0000000000000000", 15293 => "0000000000000000", 15294 => "0000000000000000", 15295 => "0000000000000000", 15296 => "0000000000000000", 15297 => "0000000000000000", 15298 => "0000000000000000", 15299 => "0000000000000000", 15300 => "0000000000000000", 15301 => "0000000000000000", 15302 => "0000000000000000", 15303 => "0000000000000000", 15304 => "0000000000000000", 15305 => "0000000000000000", 15306 => "0000000000000000", 15307 => "0000000000000000", 15308 => "0000000000000000", 15309 => "0000000000000000", 15310 => "0000000000000000", 15311 => "0000000000000000", 15312 => "0000000000000000", 15313 => "0000000000000000", 15314 => "0000000000000000", 15315 => "0000000000000000", 15316 => "0000000000000000", 15317 => "0000000000000000", 15318 => "0000000000000000", 15319 => "0000000000000000", 15320 => "0000000000000000", 15321 => "0000000000000000", 15322 => "0000000000000000", 15323 => "0000000000000000", 15324 => "0000000000000000", 15325 => "0000000000000000", 15326 => "0000000000000000", 15327 => "0000000000000000", 15328 => "0000000000000000", 15329 => "0000000000000000", 15330 => "0000000000000000", 15331 => "0000000000000000", 15332 => "0000000000000000", 15333 => "0000000000000000", 15334 => "0000000000000000", 15335 => "0000000000000000", 15336 => "0000000000000000", 15337 => "0000000000000000", 15338 => "0000000000000000", 15339 => "0000000000000000", 15340 => "0000000000000000", 15341 => "0000000000000000", 15342 => "0000000000000000", 15343 => "0000000000000000", 15344 => "0000000000000000", 15345 => "0000000000000000", 15346 => "0000000000000000", 15347 => "0000000000000000", 15348 => "0000000000000000", 15349 => "0000000000000000", 15350 => "0000000000000000", 15351 => "0000000000000000", 15352 => "0000000000000000", 15353 => "0000000000000000", 15354 => "0000000000000000", 15355 => "0000000000000000", 15356 => "0000000000000000", 15357 => "0000000000000000", 15358 => "0000000000000000", 15359 => "0000000000000000", 15360 => "0000000000000000", 15361 => "0000000000000000", 15362 => "0000000000000000", 15363 => "0000000000000000", 15364 => "0000000000000000", 15365 => "0000000000000000", 15366 => "0000000000000000", 15367 => "0000000000000000", 15368 => "0000000000000000", 15369 => "0000000000000000", 15370 => "0000000000000000", 15371 => "0000000000000000", 15372 => "0000000000000000", 15373 => "0000000000000000", 15374 => "0000000000000000", 15375 => "0000000000000000", 15376 => "0000000000000000", 15377 => "0000000000000000", 15378 => "0000000000000000", 15379 => "0000000000000000", 15380 => "0000000000000000", 15381 => "0000000000000000", 15382 => "0000000000000000", 15383 => "0000000000000000", 15384 => "0000000000000000", 15385 => "0000000000000000", 15386 => "0000000000000000", 15387 => "0000000000000000", 15388 => "0000000000000000", 15389 => "0000000000000000", 15390 => "0000000000000000", 15391 => "0000000000000000", 15392 => "0000000000000000", 15393 => "0000000000000000", 15394 => "0000000000000000", 15395 => "0000000000000000", 15396 => "0000000000000000", 15397 => "0000000000000000", 15398 => "0000000000000000", 15399 => "0000000000000000", 15400 => "0000000000000000", 15401 => "0000000000000000", 15402 => "0000000000000000", 15403 => "0000000000000000", 15404 => "0000000000000000", 15405 => "0000000000000000", 15406 => "0000000000000000", 15407 => "0000000000000000", 15408 => "0000000000000000", 15409 => "0000000000000000", 15410 => "0000000000000000", 15411 => "0000000000000000", 15412 => "0000000000000000", 15413 => "0000000000000000", 15414 => "0000000000000000", 15415 => "0000000000000000", 15416 => "0000000000000000", 15417 => "0000000000000000", 15418 => "0000000000000000", 15419 => "0000000000000000", 15420 => "0000000000000000", 15421 => "0000000000000000", 15422 => "0000000000000000", 15423 => "0000000000000000", 15424 => "0000000000000000", 15425 => "0000000000000000", 15426 => "0000000000000000", 15427 => "0000000000000000", 15428 => "0000000000000000", 15429 => "0000000000000000", 15430 => "0000000000000000", 15431 => "0000000000000000", 15432 => "0000000000000000", 15433 => "0000000000000000", 15434 => "0000000000000000", 15435 => "0000000000000000", 15436 => "0000000000000000", 15437 => "0000000000000000", 15438 => "0000000000000000", 15439 => "0000000000000000", 15440 => "0000000000000000", 15441 => "0000000000000000", 15442 => "0000000000000000", 15443 => "0000000000000000", 15444 => "0000000000000000", 15445 => "0000000000000000", 15446 => "0000000000000000", 15447 => "0000000000000000", 15448 => "0000000000000000", 15449 => "0000000000000000", 15450 => "0000000000000000", 15451 => "0000000000000000", 15452 => "0000000000000000", 15453 => "0000000000000000", 15454 => "0000000000000000", 15455 => "0000000000000000", 15456 => "0000000000000000", 15457 => "0000000000000000", 15458 => "0000000000000000", 15459 => "0000000000000000", 15460 => "0000000000000000", 15461 => "0000000000000000", 15462 => "0000000000000000", 15463 => "0000000000000000", 15464 => "0000000000000000", 15465 => "0000000000000000", 15466 => "0000000000000000", 15467 => "0000000000000000", 15468 => "0000000000000000", 15469 => "0000000000000000", 15470 => "0000000000000000", 15471 => "0000000000000000", 15472 => "0000000000000000", 15473 => "0000000000000000", 15474 => "0000000000000000", 15475 => "0000000000000000", 15476 => "0000000000000000", 15477 => "0000000000000000", 15478 => "0000000000000000", 15479 => "0000000000000000", 15480 => "0000000000000000", 15481 => "0000000000000000", 15482 => "0000000000000000", 15483 => "0000000000000000", 15484 => "0000000000000000", 15485 => "0000000000000000", 15486 => "0000000000000000", 15487 => "0000000000000000", 15488 => "0000000000000000", 15489 => "0000000000000000", 15490 => "0000000000000000", 15491 => "0000000000000000", 15492 => "0000000000000000", 15493 => "0000000000000000", 15494 => "0000000000000000", 15495 => "0000000000000000", 15496 => "0000000000000000", 15497 => "0000000000000000", 15498 => "0000000000000000", 15499 => "0000000000000000", 15500 => "0000000000000000", 15501 => "0000000000000000", 15502 => "0000000000000000", 15503 => "0000000000000000", 15504 => "0000000000000000", 15505 => "0000000000000000", 15506 => "0000000000000000", 15507 => "0000000000000000", 15508 => "0000000000000000", 15509 => "0000000000000000", 15510 => "0000000000000000", 15511 => "0000000000000000", 15512 => "0000000000000000", 15513 => "0000000000000000", 15514 => "0000000000000000", 15515 => "0000000000000000", 15516 => "0000000000000000", 15517 => "0000000000000000", 15518 => "0000000000000000", 15519 => "0000000000000000", 15520 => "0000000000000000", 15521 => "0000000000000000", 15522 => "0000000000000000", 15523 => "0000000000000000", 15524 => "0000000000000000", 15525 => "0000000000000000", 15526 => "0000000000000000", 15527 => "0000000000000000", 15528 => "0000000000000000", 15529 => "0000000000000000", 15530 => "0000000000000000", 15531 => "0000000000000000", 15532 => "0000000000000000", 15533 => "0000000000000000", 15534 => "0000000000000000", 15535 => "0000000000000000", 15536 => "0000000000000000", 15537 => "0000000000000000", 15538 => "0000000000000000", 15539 => "0000000000000000", 15540 => "0000000000000000", 15541 => "0000000000000000", 15542 => "0000000000000000", 15543 => "0000000000000000", 15544 => "0000000000000000", 15545 => "0000000000000000", 15546 => "0000000000000000", 15547 => "0000000000000000", 15548 => "0000000000000000", 15549 => "0000000000000000", 15550 => "0000000000000000", 15551 => "0000000000000000", 15552 => "0000000000000000", 15553 => "0000000000000000", 15554 => "0000000000000000", 15555 => "0000000000000000", 15556 => "0000000000000000", 15557 => "0000000000000000", 15558 => "0000000000000000", 15559 => "0000000000000000", 15560 => "0000000000000000", 15561 => "0000000000000000", 15562 => "0000000000000000", 15563 => "0000000000000000", 15564 => "0000000000000000", 15565 => "0000000000000000", 15566 => "0000000000000000", 15567 => "0000000000000000", 15568 => "0000000000000000", 15569 => "0000000000000000", 15570 => "0000000000000000", 15571 => "0000000000000000", 15572 => "0000000000000000", 15573 => "0000000000000000", 15574 => "0000000000000000", 15575 => "0000000000000000", 15576 => "0000000000000000", 15577 => "0000000000000000", 15578 => "0000000000000000", 15579 => "0000000000000000", 15580 => "0000000000000000", 15581 => "0000000000000000", 15582 => "0000000000000000", 15583 => "0000000000000000", 15584 => "0000000000000000", 15585 => "0000000000000000", 15586 => "0000000000000000", 15587 => "0000000000000000", 15588 => "0000000000000000", 15589 => "0000000000000000", 15590 => "0000000000000000", 15591 => "0000000000000000", 15592 => "0000000000000000", 15593 => "0000000000000000", 15594 => "0000000000000000", 15595 => "0000000000000000", 15596 => "0000000000000000", 15597 => "0000000000000000", 15598 => "0000000000000000", 15599 => "0000000000000000", 15600 => "0000000000000000", 15601 => "0000000000000000", 15602 => "0000000000000000", 15603 => "0000000000000000", 15604 => "0000000000000000", 15605 => "0000000000000000", 15606 => "0000000000000000", 15607 => "0000000000000000", 15608 => "0000000000000000", 15609 => "0000000000000000", 15610 => "0000000000000000", 15611 => "0000000000000000", 15612 => "0000000000000000", 15613 => "0000000000000000", 15614 => "0000000000000000", 15615 => "0000000000000000", 15616 => "0000000000000000", 15617 => "0000000000000000", 15618 => "0000000000000000", 15619 => "0000000000000000", 15620 => "0000000000000000", 15621 => "0000000000000000", 15622 => "0000000000000000", 15623 => "0000000000000000", 15624 => "0000000000000000", 15625 => "0000000000000000", 15626 => "0000000000000000", 15627 => "0000000000000000", 15628 => "0000000000000000", 15629 => "0000000000000000", 15630 => "0000000000000000", 15631 => "0000000000000000", 15632 => "0000000000000000", 15633 => "0000000000000000", 15634 => "0000000000000000", 15635 => "0000000000000000", 15636 => "0000000000000000", 15637 => "0000000000000000", 15638 => "0000000000000000", 15639 => "0000000000000000", 15640 => "0000000000000000", 15641 => "0000000000000000", 15642 => "0000000000000000", 15643 => "0000000000000000", 15644 => "0000000000000000", 15645 => "0000000000000000", 15646 => "0000000000000000", 15647 => "0000000000000000", 15648 => "0000000000000000", 15649 => "0000000000000000", 15650 => "0000000000000000", 15651 => "0000000000000000", 15652 => "0000000000000000", 15653 => "0000000000000000", 15654 => "0000000000000000", 15655 => "0000000000000000", 15656 => "0000000000000000", 15657 => "0000000000000000", 15658 => "0000000000000000", 15659 => "0000000000000000", 15660 => "0000000000000000", 15661 => "0000000000000000", 15662 => "0000000000000000", 15663 => "0000000000000000", 15664 => "0000000000000000", 15665 => "0000000000000000", 15666 => "0000000000000000", 15667 => "0000000000000000", 15668 => "0000000000000000", 15669 => "0000000000000000", 15670 => "0000000000000000", 15671 => "0000000000000000", 15672 => "0000000000000000", 15673 => "0000000000000000", 15674 => "0000000000000000", 15675 => "0000000000000000", 15676 => "0000000000000000", 15677 => "0000000000000000", 15678 => "0000000000000000", 15679 => "0000000000000000", 15680 => "0000000000000000", 15681 => "0000000000000000", 15682 => "0000000000000000", 15683 => "0000000000000000", 15684 => "0000000000000000", 15685 => "0000000000000000", 15686 => "0000000000000000", 15687 => "0000000000000000", 15688 => "0000000000000000", 15689 => "0000000000000000", 15690 => "0000000000000000", 15691 => "0000000000000000", 15692 => "0000000000000000", 15693 => "0000000000000000", 15694 => "0000000000000000", 15695 => "0000000000000000", 15696 => "0000000000000000", 15697 => "0000000000000000", 15698 => "0000000000000000", 15699 => "0000000000000000", 15700 => "0000000000000000", 15701 => "0000000000000000", 15702 => "0000000000000000", 15703 => "0000000000000000", 15704 => "0000000000000000", 15705 => "0000000000000000", 15706 => "0000000000000000", 15707 => "0000000000000000", 15708 => "0000000000000000", 15709 => "0000000000000000", 15710 => "0000000000000000", 15711 => "0000000000000000", 15712 => "0000000000000000", 15713 => "0000000000000000", 15714 => "0000000000000000", 15715 => "0000000000000000", 15716 => "0000000000000000", 15717 => "0000000000000000", 15718 => "0000000000000000", 15719 => "0000000000000000", 15720 => "0000000000000000", 15721 => "0000000000000000", 15722 => "0000000000000000", 15723 => "0000000000000000", 15724 => "0000000000000000", 15725 => "0000000000000000", 15726 => "0000000000000000", 15727 => "0000000000000000", 15728 => "0000000000000000", 15729 => "0000000000000000", 15730 => "0000000000000000", 15731 => "0000000000000000", 15732 => "0000000000000000", 15733 => "0000000000000000", 15734 => "0000000000000000", 15735 => "0000000000000000", 15736 => "0000000000000000", 15737 => "0000000000000000", 15738 => "0000000000000000", 15739 => "0000000000000000", 15740 => "0000000000000000", 15741 => "0000000000000000", 15742 => "0000000000000000", 15743 => "0000000000000000", 15744 => "0000000000000000", 15745 => "0000000000000000", 15746 => "0000000000000000", 15747 => "0000000000000000", 15748 => "0000000000000000", 15749 => "0000000000000000", 15750 => "0000000000000000", 15751 => "0000000000000000", 15752 => "0000000000000000", 15753 => "0000000000000000", 15754 => "0000000000000000", 15755 => "0000000000000000", 15756 => "0000000000000000", 15757 => "0000000000000000", 15758 => "0000000000000000", 15759 => "0000000000000000", 15760 => "0000000000000000", 15761 => "0000000000000000", 15762 => "0000000000000000", 15763 => "0000000000000000", 15764 => "0000000000000000", 15765 => "0000000000000000", 15766 => "0000000000000000", 15767 => "0000000000000000", 15768 => "0000000000000000", 15769 => "0000000000000000", 15770 => "0000000000000000", 15771 => "0000000000000000", 15772 => "0000000000000000", 15773 => "0000000000000000", 15774 => "0000000000000000", 15775 => "0000000000000000", 15776 => "0000000000000000", 15777 => "0000000000000000", 15778 => "0000000000000000", 15779 => "0000000000000000", 15780 => "0000000000000000", 15781 => "0000000000000000", 15782 => "0000000000000000", 15783 => "0000000000000000", 15784 => "0000000000000000", 15785 => "0000000000000000", 15786 => "0000000000000000", 15787 => "0000000000000000", 15788 => "0000000000000000", 15789 => "0000000000000000", 15790 => "0000000000000000", 15791 => "0000000000000000", 15792 => "0000000000000000", 15793 => "0000000000000000", 15794 => "0000000000000000", 15795 => "0000000000000000", 15796 => "0000000000000000", 15797 => "0000000000000000", 15798 => "0000000000000000", 15799 => "0000000000000000", 15800 => "0000000000000000", 15801 => "0000000000000000", 15802 => "0000000000000000", 15803 => "0000000000000000", 15804 => "0000000000000000", 15805 => "0000000000000000", 15806 => "0000000000000000", 15807 => "0000000000000000", 15808 => "0000000000000000", 15809 => "0000000000000000", 15810 => "0000000000000000", 15811 => "0000000000000000", 15812 => "0000000000000000", 15813 => "0000000000000000", 15814 => "0000000000000000", 15815 => "0000000000000000", 15816 => "0000000000000000", 15817 => "0000000000000000", 15818 => "0000000000000000", 15819 => "0000000000000000", 15820 => "0000000000000000", 15821 => "0000000000000000", 15822 => "0000000000000000", 15823 => "0000000000000000", 15824 => "0000000000000000", 15825 => "0000000000000000", 15826 => "0000000000000000", 15827 => "0000000000000000", 15828 => "0000000000000000", 15829 => "0000000000000000", 15830 => "0000000000000000", 15831 => "0000000000000000", 15832 => "0000000000000000", 15833 => "0000000000000000", 15834 => "0000000000000000", 15835 => "0000000000000000", 15836 => "0000000000000000", 15837 => "0000000000000000", 15838 => "0000000000000000", 15839 => "0000000000000000", 15840 => "0000000000000000", 15841 => "0000000000000000", 15842 => "0000000000000000", 15843 => "0000000000000000", 15844 => "0000000000000000", 15845 => "0000000000000000", 15846 => "0000000000000000", 15847 => "0000000000000000", 15848 => "0000000000000000", 15849 => "0000000000000000", 15850 => "0000000000000000", 15851 => "0000000000000000", 15852 => "0000000000000000", 15853 => "0000000000000000", 15854 => "0000000000000000", 15855 => "0000000000000000", 15856 => "0000000000000000", 15857 => "0000000000000000", 15858 => "0000000000000000", 15859 => "0000000000000000", 15860 => "0000000000000000", 15861 => "0000000000000000", 15862 => "0000000000000000", 15863 => "0000000000000000", 15864 => "0000000000000000", 15865 => "0000000000000000", 15866 => "0000000000000000", 15867 => "0000000000000000", 15868 => "0000000000000000", 15869 => "0000000000000000", 15870 => "0000000000000000", 15871 => "0000000000000000", 15872 => "0000000000000000", 15873 => "0000000000000000", 15874 => "0000000000000000", 15875 => "0000000000000000", 15876 => "0000000000000000", 15877 => "0000000000000000", 15878 => "0000000000000000", 15879 => "0000000000000000", 15880 => "0000000000000000", 15881 => "0000000000000000", 15882 => "0000000000000000", 15883 => "0000000000000000", 15884 => "0000000000000000", 15885 => "0000000000000000", 15886 => "0000000000000000", 15887 => "0000000000000000", 15888 => "0000000000000000", 15889 => "0000000000000000", 15890 => "0000000000000000", 15891 => "0000000000000000", 15892 => "0000000000000000", 15893 => "0000000000000000", 15894 => "0000000000000000", 15895 => "0000000000000000", 15896 => "0000000000000000", 15897 => "0000000000000000", 15898 => "0000000000000000", 15899 => "0000000000000000", 15900 => "0000000000000000", 15901 => "0000000000000000", 15902 => "0000000000000000", 15903 => "0000000000000000", 15904 => "0000000000000000", 15905 => "0000000000000000", 15906 => "0000000000000000", 15907 => "0000000000000000", 15908 => "0000000000000000", 15909 => "0000000000000000", 15910 => "0000000000000000", 15911 => "0000000000000000", 15912 => "0000000000000000", 15913 => "0000000000000000", 15914 => "0000000000000000", 15915 => "0000000000000000", 15916 => "0000000000000000", 15917 => "0000000000000000", 15918 => "0000000000000000", 15919 => "0000000000000000", 15920 => "0000000000000000", 15921 => "0000000000000000", 15922 => "0000000000000000", 15923 => "0000000000000000", 15924 => "0000000000000000", 15925 => "0000000000000000", 15926 => "0000000000000000", 15927 => "0000000000000000", 15928 => "0000000000000000", 15929 => "0000000000000000", 15930 => "0000000000000000", 15931 => "0000000000000000", 15932 => "0000000000000000", 15933 => "0000000000000000", 15934 => "0000000000000000", 15935 => "0000000000000000", 15936 => "0000000000000000", 15937 => "0000000000000000", 15938 => "0000000000000000", 15939 => "0000000000000000", 15940 => "0000000000000000", 15941 => "0000000000000000", 15942 => "0000000000000000", 15943 => "0000000000000000", 15944 => "0000000000000000", 15945 => "0000000000000000", 15946 => "0000000000000000", 15947 => "0000000000000000", 15948 => "0000000000000000", 15949 => "0000000000000000", 15950 => "0000000000000000", 15951 => "0000000000000000", 15952 => "0000000000000000", 15953 => "0000000000000000", 15954 => "0000000000000000", 15955 => "0000000000000000", 15956 => "0000000000000000", 15957 => "0000000000000000", 15958 => "0000000000000000", 15959 => "0000000000000000", 15960 => "0000000000000000", 15961 => "0000000000000000", 15962 => "0000000000000000", 15963 => "0000000000000000", 15964 => "0000000000000000", 15965 => "0000000000000000", 15966 => "0000000000000000", 15967 => "0000000000000000", 15968 => "0000000000000000", 15969 => "0000000000000000", 15970 => "0000000000000000", 15971 => "0000000000000000", 15972 => "0000000000000000", 15973 => "0000000000000000", 15974 => "0000000000000000", 15975 => "0000000000000000", 15976 => "0000000000000000", 15977 => "0000000000000000", 15978 => "0000000000000000", 15979 => "0000000000000000", 15980 => "0000000000000000", 15981 => "0000000000000000", 15982 => "0000000000000000", 15983 => "0000000000000000", 15984 => "0000000000000000", 15985 => "0000000000000000", 15986 => "0000000000000000", 15987 => "0000000000000000", 15988 => "0000000000000000", 15989 => "0000000000000000", 15990 => "0000000000000000", 15991 => "0000000000000000", 15992 => "0000000000000000", 15993 => "0000000000000000", 15994 => "0000000000000000", 15995 => "0000000000000000", 15996 => "0000000000000000", 15997 => "0000000000000000", 15998 => "0000000000000000", 15999 => "0000000000000000", 16000 => "0000000000000000", 16001 => "0000000000000000", 16002 => "0000000000000000", 16003 => "0000000000000000", 16004 => "0000000000000000", 16005 => "0000000000000000", 16006 => "0000000000000000", 16007 => "0000000000000000", 16008 => "0000000000000000", 16009 => "0000000000000000", 16010 => "0000000000000000", 16011 => "0000000000000000", 16012 => "0000000000000000", 16013 => "0000000000000000", 16014 => "0000000000000000", 16015 => "0000000000000000", 16016 => "0000000000000000", 16017 => "0000000000000000", 16018 => "0000000000000000", 16019 => "0000000000000000", 16020 => "0000000000000000", 16021 => "0000000000000000", 16022 => "0000000000000000", 16023 => "0000000000000000", 16024 => "0000000000000000", 16025 => "0000000000000000", 16026 => "0000000000000000", 16027 => "0000000000000000", 16028 => "0000000000000000", 16029 => "0000000000000000", 16030 => "0000000000000000", 16031 => "0000000000000000", 16032 => "0000000000000000", 16033 => "0000000000000000", 16034 => "0000000000000000", 16035 => "0000000000000000", 16036 => "0000000000000000", 16037 => "0000000000000000", 16038 => "0000000000000000", 16039 => "0000000000000000", 16040 => "0000000000000000", 16041 => "0000000000000000", 16042 => "0000000000000000", 16043 => "0000000000000000", 16044 => "0000000000000000", 16045 => "0000000000000000", 16046 => "0000000000000000", 16047 => "0000000000000000", 16048 => "0000000000000000", 16049 => "0000000000000000", 16050 => "0000000000000000", 16051 => "0000000000000000", 16052 => "0000000000000000", 16053 => "0000000000000000", 16054 => "0000000000000000", 16055 => "0000000000000000", 16056 => "0000000000000000", 16057 => "0000000000000000", 16058 => "0000000000000000", 16059 => "0000000000000000", 16060 => "0000000000000000", 16061 => "0000000000000000", 16062 => "0000000000000000", 16063 => "0000000000000000", 16064 => "0000000000000000", 16065 => "0000000000000000", 16066 => "0000000000000000", 16067 => "0000000000000000", 16068 => "0000000000000000", 16069 => "0000000000000000", 16070 => "0000000000000000", 16071 => "0000000000000000", 16072 => "0000000000000000", 16073 => "0000000000000000", 16074 => "0000000000000000", 16075 => "0000000000000000", 16076 => "0000000000000000", 16077 => "0000000000000000", 16078 => "0000000000000000", 16079 => "0000000000000000", 16080 => "0000000000000000", 16081 => "0000000000000000", 16082 => "0000000000000000", 16083 => "0000000000000000", 16084 => "0000000000000000", 16085 => "0000000000000000", 16086 => "0000000000000000", 16087 => "0000000000000000", 16088 => "0000000000000000", 16089 => "0000000000000000", 16090 => "0000000000000000", 16091 => "0000000000000000", 16092 => "0000000000000000", 16093 => "0000000000000000", 16094 => "0000000000000000", 16095 => "0000000000000000", 16096 => "0000000000000000", 16097 => "0000000000000000", 16098 => "0000000000000000", 16099 => "0000000000000000", 16100 => "0000000000000000", 16101 => "0000000000000000", 16102 => "0000000000000000", 16103 => "0000000000000000", 16104 => "0000000000000000", 16105 => "0000000000000000", 16106 => "0000000000000000", 16107 => "0000000000000000", 16108 => "0000000000000000", 16109 => "0000000000000000", 16110 => "0000000000000000", 16111 => "0000000000000000", 16112 => "0000000000000000", 16113 => "0000000000000000", 16114 => "0000000000000000", 16115 => "0000000000000000", 16116 => "0000000000000000", 16117 => "0000000000000000", 16118 => "0000000000000000", 16119 => "0000000000000000", 16120 => "0000000000000000", 16121 => "0000000000000000", 16122 => "0000000000000000", 16123 => "0000000000000000", 16124 => "0000000000000000", 16125 => "0000000000000000", 16126 => "0000000000000000", 16127 => "0000000000000000", 16128 => "0000000000000000", 16129 => "0000000000000000", 16130 => "0000000000000000", 16131 => "0000000000000000", 16132 => "0000000000000000", 16133 => "0000000000000000", 16134 => "0000000000000000", 16135 => "0000000000000000", 16136 => "0000000000000000", 16137 => "0000000000000000", 16138 => "0000000000000000", 16139 => "0000000000000000", 16140 => "0000000000000000", 16141 => "0000000000000000", 16142 => "0000000000000000", 16143 => "0000000000000000", 16144 => "0000000000000000", 16145 => "0000000000000000", 16146 => "0000000000000000", 16147 => "0000000000000000", 16148 => "0000000000000000", 16149 => "0000000000000000", 16150 => "0000000000000000", 16151 => "0000000000000000", 16152 => "0000000000000000", 16153 => "0000000000000000", 16154 => "0000000000000000", 16155 => "0000000000000000", 16156 => "0000000000000000", 16157 => "0000000000000000", 16158 => "0000000000000000", 16159 => "0000000000000000", 16160 => "0000000000000000", 16161 => "0000000000000000", 16162 => "0000000000000000", 16163 => "0000000000000000", 16164 => "0000000000000000", 16165 => "0000000000000000", 16166 => "0000000000000000", 16167 => "0000000000000000", 16168 => "0000000000000000", 16169 => "0000000000000000", 16170 => "0000000000000000", 16171 => "0000000000000000", 16172 => "0000000000000000", 16173 => "0000000000000000", 16174 => "0000000000000000", 16175 => "0000000000000000", 16176 => "0000000000000000", 16177 => "0000000000000000", 16178 => "0000000000000000", 16179 => "0000000000000000", 16180 => "0000000000000000", 16181 => "0000000000000000", 16182 => "0000000000000000", 16183 => "0000000000000000", 16184 => "0000000000000000", 16185 => "0000000000000000", 16186 => "0000000000000000", 16187 => "0000000000000000", 16188 => "0000000000000000", 16189 => "0000000000000000", 16190 => "0000000000000000", 16191 => "0000000000000000", 16192 => "0000000000000000", 16193 => "0000000000000000", 16194 => "0000000000000000", 16195 => "0000000000000000", 16196 => "0000000000000000", 16197 => "0000000000000000", 16198 => "0000000000000000", 16199 => "0000000000000000", 16200 => "0000000000000000", 16201 => "0000000000000000", 16202 => "0000000000000000", 16203 => "0000000000000000", 16204 => "0000000000000000", 16205 => "0000000000000000", 16206 => "0000000000000000", 16207 => "0000000000000000", 16208 => "0000000000000000", 16209 => "0000000000000000", 16210 => "0000000000000000", 16211 => "0000000000000000", 16212 => "0000000000000000", 16213 => "0000000000000000", 16214 => "0000000000000000", 16215 => "0000000000000000", 16216 => "0000000000000000", 16217 => "0000000000000000", 16218 => "0000000000000000", 16219 => "0000000000000000", 16220 => "0000000000000000", 16221 => "0000000000000000", 16222 => "0000000000000000", 16223 => "0000000000000000", 16224 => "0000000000000000", 16225 => "0000000000000000", 16226 => "0000000000000000", 16227 => "0000000000000000", 16228 => "0000000000000000", 16229 => "0000000000000000", 16230 => "0000000000000000", 16231 => "0000000000000000", 16232 => "0000000000000000", 16233 => "0000000000000000", 16234 => "0000000000000000", 16235 => "0000000000000000", 16236 => "0000000000000000", 16237 => "0000000000000000", 16238 => "0000000000000000", 16239 => "0000000000000000", 16240 => "0000000000000000", 16241 => "0000000000000000", 16242 => "0000000000000000", 16243 => "0000000000000000", 16244 => "0000000000000000", 16245 => "0000000000000000", 16246 => "0000000000000000", 16247 => "0000000000000000", 16248 => "0000000000000000", 16249 => "0000000000000000", 16250 => "0000000000000000", 16251 => "0000000000000000", 16252 => "0000000000000000", 16253 => "0000000000000000", 16254 => "0000000000000000", 16255 => "0000000000000000", 16256 => "0000000000000000", 16257 => "0000000000000000", 16258 => "0000000000000000", 16259 => "0000000000000000", 16260 => "0000000000000000", 16261 => "0000000000000000", 16262 => "0000000000000000", 16263 => "0000000000000000", 16264 => "0000000000000000", 16265 => "0000000000000000", 16266 => "0000000000000000", 16267 => "0000000000000000", 16268 => "0000000000000000", 16269 => "0000000000000000", 16270 => "0000000000000000", 16271 => "0000000000000000", 16272 => "0000000000000000", 16273 => "0000000000000000", 16274 => "0000000000000000", 16275 => "0000000000000000", 16276 => "0000000000000000", 16277 => "0000000000000000", 16278 => "0000000000000000", 16279 => "0000000000000000", 16280 => "0000000000000000", 16281 => "0000000000000000", 16282 => "0000000000000000", 16283 => "0000000000000000", 16284 => "0000000000000000", 16285 => "0000000000000000", 16286 => "0000000000000000", 16287 => "0000000000000000", 16288 => "0000000000000000", 16289 => "0000000000000000", 16290 => "0000000000000000", 16291 => "0000000000000000", 16292 => "0000000000000000", 16293 => "0000000000000000", 16294 => "0000000000000000", 16295 => "0000000000000000", 16296 => "0000000000000000", 16297 => "0000000000000000", 16298 => "0000000000000000", 16299 => "0000000000000000", 16300 => "0000000000000000", 16301 => "0000000000000000", 16302 => "0000000000000000", 16303 => "0000000000000000", 16304 => "0000000000000000", 16305 => "0000000000000000", 16306 => "0000000000000000", 16307 => "0000000000000000", 16308 => "0000000000000000", 16309 => "0000000000000000", 16310 => "0000000000000000", 16311 => "0000000000000000", 16312 => "0000000000000000", 16313 => "0000000000000000", 16314 => "0000000000000000", 16315 => "0000000000000000", 16316 => "0000000000000000", 16317 => "0000000000000000", 16318 => "0000000000000000", 16319 => "0000000000000000", 16320 => "0000000000000000", 16321 => "0000000000000000", 16322 => "0000000000000000", 16323 => "0000000000000000", 16324 => "0000000000000000", 16325 => "0000000000000000", 16326 => "0000000000000000", 16327 => "0000000000000000", 16328 => "0000000000000000", 16329 => "0000000000000000", 16330 => "0000000000000000", 16331 => "0000000000000000", 16332 => "0000000000000000", 16333 => "0000000000000000", 16334 => "0000000000000000", 16335 => "0000000000000000", 16336 => "0000000000000000", 16337 => "0000000000000000", 16338 => "0000000000000000", 16339 => "0000000000000000", 16340 => "0000000000000000", 16341 => "0000000000000000", 16342 => "0000000000000000", 16343 => "0000000000000000", 16344 => "0000000000000000", 16345 => "0000000000000000", 16346 => "0000000000000000", 16347 => "0000000000000000", 16348 => "0000000000000000", 16349 => "0000000000000000", 16350 => "0000000000000000", 16351 => "0000000000000000", 16352 => "0000000000000000", 16353 => "0000000000000000", 16354 => "0000000000000000", 16355 => "0000000000000000", 16356 => "0000000000000000", 16357 => "0000000000000000", 16358 => "0000000000000000", 16359 => "0000000000000000", 16360 => "0000000000000000", 16361 => "0000000000000000", 16362 => "0000000000000000", 16363 => "0000000000000000", 16364 => "0000000000000000", 16365 => "0000000000000000", 16366 => "0000000000000000", 16367 => "0000000000000000", 16368 => "0000000000000000", 16369 => "0000000000000000", 16370 => "0000000000000000", 16371 => "0000000000000000", 16372 => "0000000000000000", 16373 => "0000000000000000", 16374 => "0000000000000000", 16375 => "0000000000000000", 16376 => "0000000000000000", 16377 => "0000000000000000", 16378 => "0000000000000000", 16379 => "0000000000000000", 16380 => "0000000000000000", 16381 => "0000000000000000", 16382 => "0000000000000000", 16383 => "0000000000000000", 16384 => "0000000000000000", 16385 => "0000000000000000", 16386 => "0000000000000000", 16387 => "0000000000000000", 16388 => "0000000000000000", 16389 => "0000000000000000", 16390 => "0000000000000000", 16391 => "0000000000000000", 16392 => "0000000000000000", 16393 => "0000000000000000", 16394 => "0000000000000000", 16395 => "0000000000000000", 16396 => "0000000000000000", 16397 => "0000000000000000", 16398 => "0000000000000000", 16399 => "0000000000000000", 16400 => "0000000000000000", 16401 => "0000000000000000", 16402 => "0000000000000000", 16403 => "0000000000000000", 16404 => "0000000000000000", 16405 => "0000000000000000", 16406 => "0000000000000000", 16407 => "0000000000000000", 16408 => "0000000000000000", 16409 => "0000000000000000", 16410 => "0000000000000000", 16411 => "0000000000000000", 16412 => "0000000000000000", 16413 => "0000000000000000", 16414 => "0000000000000000", 16415 => "0000000000000000", 16416 => "0000000000000000", 16417 => "0000000000000000", 16418 => "0000000000000000", 16419 => "0000000000000000", 16420 => "0000000000000000", 16421 => "0000000000000000", 16422 => "0000000000000000", 16423 => "0000000000000000", 16424 => "0000000000000000", 16425 => "0000000000000000", 16426 => "0000000000000000", 16427 => "0000000000000000", 16428 => "0000000000000000", 16429 => "0000000000000000", 16430 => "0000000000000000", 16431 => "0000000000000000", 16432 => "0000000000000000", 16433 => "0000000000000000", 16434 => "0000000000000000", 16435 => "0000000000000000", 16436 => "0000000000000000", 16437 => "0000000000000000", 16438 => "0000000000000000", 16439 => "0000000000000000", 16440 => "0000000000000000", 16441 => "0000000000000000", 16442 => "0000000000000000", 16443 => "0000000000000000", 16444 => "0000000000000000", 16445 => "0000000000000000", 16446 => "0000000000000000", 16447 => "0000000000000000", 16448 => "0000000000000000", 16449 => "0000000000000000", 16450 => "0000000000000000", 16451 => "0000000000000000", 16452 => "0000000000000000", 16453 => "0000000000000000", 16454 => "0000000000000000", 16455 => "0000000000000000", 16456 => "0000000000000000", 16457 => "0000000000000000", 16458 => "0000000000000000", 16459 => "0000000000000000", 16460 => "0000000000000000", 16461 => "0000000000000000", 16462 => "0000000000000000", 16463 => "0000000000000000", 16464 => "0000000000000000", 16465 => "0000000000000000", 16466 => "0000000000000000", 16467 => "0000000000000000", 16468 => "0000000000000000", 16469 => "0000000000000000", 16470 => "0000000000000000", 16471 => "0000000000000000", 16472 => "0000000000000000", 16473 => "0000000000000000", 16474 => "0000000000000000", 16475 => "0000000000000000", 16476 => "0000000000000000", 16477 => "0000000000000000", 16478 => "0000000000000000", 16479 => "0000000000000000", 16480 => "0000000000000000", 16481 => "0000000000000000", 16482 => "0000000000000000", 16483 => "0000000000000000", 16484 => "0000000000000000", 16485 => "0000000000000000", 16486 => "0000000000000000", 16487 => "0000000000000000", 16488 => "0000000000000000", 16489 => "0000000000000000", 16490 => "0000000000000000", 16491 => "0000000000000000", 16492 => "0000000000000000", 16493 => "0000000000000000", 16494 => "0000000000000000", 16495 => "0000000000000000", 16496 => "0000000000000000", 16497 => "0000000000000000", 16498 => "0000000000000000", 16499 => "0000000000000000", 16500 => "0000000000000000", 16501 => "0000000000000000", 16502 => "0000000000000000", 16503 => "0000000000000000", 16504 => "0000000000000000", 16505 => "0000000000000000", 16506 => "0000000000000000", 16507 => "0000000000000000", 16508 => "0000000000000000", 16509 => "0000000000000000", 16510 => "0000000000000000", 16511 => "0000000000000000", 16512 => "0000000000000000", 16513 => "0000000000000000", 16514 => "0000000000000000", 16515 => "0000000000000000", 16516 => "0000000000000000", 16517 => "0000000000000000", 16518 => "0000000000000000", 16519 => "0000000000000000", 16520 => "0000000000000000", 16521 => "0000000000000000", 16522 => "0000000000000000", 16523 => "0000000000000000", 16524 => "0000000000000000", 16525 => "0000000000000000", 16526 => "0000000000000000", 16527 => "0000000000000000", 16528 => "0000000000000000", 16529 => "0000000000000000", 16530 => "0000000000000000", 16531 => "0000000000000000", 16532 => "0000000000000000", 16533 => "0000000000000000", 16534 => "0000000000000000", 16535 => "0000000000000000", 16536 => "0000000000000000", 16537 => "0000000000000000", 16538 => "0000000000000000", 16539 => "0000000000000000", 16540 => "0000000000000000", 16541 => "0000000000000000", 16542 => "0000000000000000", 16543 => "0000000000000000", 16544 => "0000000000000000", 16545 => "0000000000000000", 16546 => "0000000000000000", 16547 => "0000000000000000", 16548 => "0000000000000000", 16549 => "0000000000000000", 16550 => "0000000000000000", 16551 => "0000000000000000", 16552 => "0000000000000000", 16553 => "0000000000000000", 16554 => "0000000000000000", 16555 => "0000000000000000", 16556 => "0000000000000000", 16557 => "0000000000000000", 16558 => "0000000000000000", 16559 => "0000000000000000", 16560 => "0000000000000000", 16561 => "0000000000000000", 16562 => "0000000000000000", 16563 => "0000000000000000", 16564 => "0000000000000000", 16565 => "0000000000000000", 16566 => "0000000000000000", 16567 => "0000000000000000", 16568 => "0000000000000000", 16569 => "0000000000000000", 16570 => "0000000000000000", 16571 => "0000000000000000", 16572 => "0000000000000000", 16573 => "0000000000000000", 16574 => "0000000000000000", 16575 => "0000000000000000", 16576 => "0000000000000000", 16577 => "0000000000000000", 16578 => "0000000000000000", 16579 => "0000000000000000", 16580 => "0000000000000000", 16581 => "0000000000000000", 16582 => "0000000000000000", 16583 => "0000000000000000", 16584 => "0000000000000000", 16585 => "0000000000000000", 16586 => "0000000000000000", 16587 => "0000000000000000", 16588 => "0000000000000000", 16589 => "0000000000000000", 16590 => "0000000000000000", 16591 => "0000000000000000", 16592 => "0000000000000000", 16593 => "0000000000000000", 16594 => "0000000000000000", 16595 => "0000000000000000", 16596 => "0000000000000000", 16597 => "0000000000000000", 16598 => "0000000000000000", 16599 => "0000000000000000", 16600 => "0000000000000000", 16601 => "0000000000000000", 16602 => "0000000000000000", 16603 => "0000000000000000", 16604 => "0000000000000000", 16605 => "0000000000000000", 16606 => "0000000000000000", 16607 => "0000000000000000", 16608 => "0000000000000000", 16609 => "0000000000000000", 16610 => "0000000000000000", 16611 => "0000000000000000", 16612 => "0000000000000000", 16613 => "0000000000000000", 16614 => "0000000000000000", 16615 => "0000000000000000", 16616 => "0000000000000000", 16617 => "0000000000000000", 16618 => "0000000000000000", 16619 => "0000000000000000", 16620 => "0000000000000000", 16621 => "0000000000000000", 16622 => "0000000000000000", 16623 => "0000000000000000", 16624 => "0000000000000000", 16625 => "0000000000000000", 16626 => "0000000000000000", 16627 => "0000000000000000", 16628 => "0000000000000000", 16629 => "0000000000000000", 16630 => "0000000000000000", 16631 => "0000000000000000", 16632 => "0000000000000000", 16633 => "0000000000000000", 16634 => "0000000000000000", 16635 => "0000000000000000", 16636 => "0000000000000000", 16637 => "0000000000000000", 16638 => "0000000000000000", 16639 => "0000000000000000", 16640 => "0000000000000000", 16641 => "0000000000000000", 16642 => "0000000000000000", 16643 => "0000000000000000", 16644 => "0000000000000000", 16645 => "0000000000000000", 16646 => "0000000000000000", 16647 => "0000000000000000", 16648 => "0000000000000000", 16649 => "0000000000000000", 16650 => "0000000000000000", 16651 => "0000000000000000", 16652 => "0000000000000000", 16653 => "0000000000000000", 16654 => "0000000000000000", 16655 => "0000000000000000", 16656 => "0000000000000000", 16657 => "0000000000000000", 16658 => "0000000000000000", 16659 => "0000000000000000", 16660 => "0000000000000000", 16661 => "0000000000000000", 16662 => "0000000000000000", 16663 => "0000000000000000", 16664 => "0000000000000000", 16665 => "0000000000000000", 16666 => "0000000000000000", 16667 => "0000000000000000", 16668 => "0000000000000000", 16669 => "0000000000000000", 16670 => "0000000000000000", 16671 => "0000000000000000", 16672 => "0000000000000000", 16673 => "0000000000000000", 16674 => "0000000000000000", 16675 => "0000000000000000", 16676 => "0000000000000000", 16677 => "0000000000000000", 16678 => "0000000000000000", 16679 => "0000000000000000", 16680 => "0000000000000000", 16681 => "0000000000000000", 16682 => "0000000000000000", 16683 => "0000000000000000", 16684 => "0000000000000000", 16685 => "0000000000000000", 16686 => "0000000000000000", 16687 => "0000000000000000", 16688 => "0000000000000000", 16689 => "0000000000000000", 16690 => "0000000000000000", 16691 => "0000000000000000", 16692 => "0000000000000000", 16693 => "0000000000000000", 16694 => "0000000000000000", 16695 => "0000000000000000", 16696 => "0000000000000000", 16697 => "0000000000000000", 16698 => "0000000000000000", 16699 => "0000000000000000", 16700 => "0000000000000000", 16701 => "0000000000000000", 16702 => "0000000000000000", 16703 => "0000000000000000", 16704 => "0000000000000000", 16705 => "0000000000000000", 16706 => "0000000000000000", 16707 => "0000000000000000", 16708 => "0000000000000000", 16709 => "0000000000000000", 16710 => "0000000000000000", 16711 => "0000000000000000", 16712 => "0000000000000000", 16713 => "0000000000000000", 16714 => "0000000000000000", 16715 => "0000000000000000", 16716 => "0000000000000000", 16717 => "0000000000000000", 16718 => "0000000000000000", 16719 => "0000000000000000", 16720 => "0000000000000000", 16721 => "0000000000000000", 16722 => "0000000000000000", 16723 => "0000000000000000", 16724 => "0000000000000000", 16725 => "0000000000000000", 16726 => "0000000000000000", 16727 => "0000000000000000", 16728 => "0000000000000000", 16729 => "0000000000000000", 16730 => "0000000000000000", 16731 => "0000000000000000", 16732 => "0000000000000000", 16733 => "0000000000000000", 16734 => "0000000000000000", 16735 => "0000000000000000", 16736 => "0000000000000000", 16737 => "0000000000000000", 16738 => "0000000000000000", 16739 => "0000000000000000", 16740 => "0000000000000000", 16741 => "0000000000000000", 16742 => "0000000000000000", 16743 => "0000000000000000", 16744 => "0000000000000000", 16745 => "0000000000000000", 16746 => "0000000000000000", 16747 => "0000000000000000", 16748 => "0000000000000000", 16749 => "0000000000000000", 16750 => "0000000000000000", 16751 => "0000000000000000", 16752 => "0000000000000000", 16753 => "0000000000000000", 16754 => "0000000000000000", 16755 => "0000000000000000", 16756 => "0000000000000000", 16757 => "0000000000000000", 16758 => "0000000000000000", 16759 => "0000000000000000", 16760 => "0000000000000000", 16761 => "0000000000000000", 16762 => "0000000000000000", 16763 => "0000000000000000", 16764 => "0000000000000000", 16765 => "0000000000000000", 16766 => "0000000000000000", 16767 => "0000000000000000", 16768 => "0000000000000000", 16769 => "0000000000000000", 16770 => "0000000000000000", 16771 => "0000000000000000", 16772 => "0000000000000000", 16773 => "0000000000000000", 16774 => "0000000000000000", 16775 => "0000000000000000", 16776 => "0000000000000000", 16777 => "0000000000000000", 16778 => "0000000000000000", 16779 => "0000000000000000", 16780 => "0000000000000000", 16781 => "0000000000000000", 16782 => "0000000000000000", 16783 => "0000000000000000", 16784 => "0000000000000000", 16785 => "0000000000000000", 16786 => "0000000000000000", 16787 => "0000000000000000", 16788 => "0000000000000000", 16789 => "0000000000000000", 16790 => "0000000000000000", 16791 => "0000000000000000", 16792 => "0000000000000000", 16793 => "0000000000000000", 16794 => "0000000000000000", 16795 => "0000000000000000", 16796 => "0000000000000000", 16797 => "0000000000000000", 16798 => "0000000000000000", 16799 => "0000000000000000", 16800 => "0000000000000000", 16801 => "0000000000000000", 16802 => "0000000000000000", 16803 => "0000000000000000", 16804 => "0000000000000000", 16805 => "0000000000000000", 16806 => "0000000000000000", 16807 => "0000000000000000", 16808 => "0000000000000000", 16809 => "0000000000000000", 16810 => "0000000000000000", 16811 => "0000000000000000", 16812 => "0000000000000000", 16813 => "0000000000000000", 16814 => "0000000000000000", 16815 => "0000000000000000", 16816 => "0000000000000000", 16817 => "0000000000000000", 16818 => "0000000000000000", 16819 => "0000000000000000", 16820 => "0000000000000000", 16821 => "0000000000000000", 16822 => "0000000000000000", 16823 => "0000000000000000", 16824 => "0000000000000000", 16825 => "0000000000000000", 16826 => "0000000000000000", 16827 => "0000000000000000", 16828 => "0000000000000000", 16829 => "0000000000000000", 16830 => "0000000000000000", 16831 => "0000000000000000", 16832 => "0000000000000000", 16833 => "0000000000000000", 16834 => "0000000000000000", 16835 => "0000000000000000", 16836 => "0000000000000000", 16837 => "0000000000000000", 16838 => "0000000000000000", 16839 => "0000000000000000", 16840 => "0000000000000000", 16841 => "0000000000000000", 16842 => "0000000000000000", 16843 => "0000000000000000", 16844 => "0000000000000000", 16845 => "0000000000000000", 16846 => "0000000000000000", 16847 => "0000000000000000", 16848 => "0000000000000000", 16849 => "0000000000000000", 16850 => "0000000000000000", 16851 => "0000000000000000", 16852 => "0000000000000000", 16853 => "0000000000000000", 16854 => "0000000000000000", 16855 => "0000000000000000", 16856 => "0000000000000000", 16857 => "0000000000000000", 16858 => "0000000000000000", 16859 => "0000000000000000", 16860 => "0000000000000000", 16861 => "0000000000000000", 16862 => "0000000000000000", 16863 => "0000000000000000", 16864 => "0000000000000000", 16865 => "0000000000000000", 16866 => "0000000000000000", 16867 => "0000000000000000", 16868 => "0000000000000000", 16869 => "0000000000000000", 16870 => "0000000000000000", 16871 => "0000000000000000", 16872 => "0000000000000000", 16873 => "0000000000000000", 16874 => "0000000000000000", 16875 => "0000000000000000", 16876 => "0000000000000000", 16877 => "0000000000000000", 16878 => "0000000000000000", 16879 => "0000000000000000", 16880 => "0000000000000000", 16881 => "0000000000000000", 16882 => "0000000000000000", 16883 => "0000000000000000", 16884 => "0000000000000000", 16885 => "0000000000000000", 16886 => "0000000000000000", 16887 => "0000000000000000", 16888 => "0000000000000000", 16889 => "0000000000000000", 16890 => "0000000000000000", 16891 => "0000000000000000", 16892 => "0000000000000000", 16893 => "0000000000000000", 16894 => "0000000000000000", 16895 => "0000000000000000", 16896 => "0000000000000000", 16897 => "0000000000000000", 16898 => "0000000000000000", 16899 => "0000000000000000", 16900 => "0000000000000000", 16901 => "0000000000000000", 16902 => "0000000000000000", 16903 => "0000000000000000", 16904 => "0000000000000000", 16905 => "0000000000000000", 16906 => "0000000000000000", 16907 => "0000000000000000", 16908 => "0000000000000000", 16909 => "0000000000000000", 16910 => "0000000000000000", 16911 => "0000000000000000", 16912 => "0000000000000000", 16913 => "0000000000000000", 16914 => "0000000000000000", 16915 => "0000000000000000", 16916 => "0000000000000000", 16917 => "0000000000000000", 16918 => "0000000000000000", 16919 => "0000000000000000", 16920 => "0000000000000000", 16921 => "0000000000000000", 16922 => "0000000000000000", 16923 => "0000000000000000", 16924 => "0000000000000000", 16925 => "0000000000000000", 16926 => "0000000000000000", 16927 => "0000000000000000", 16928 => "0000000000000000", 16929 => "0000000000000000", 16930 => "0000000000000000", 16931 => "0000000000000000", 16932 => "0000000000000000", 16933 => "0000000000000000", 16934 => "0000000000000000", 16935 => "0000000000000000", 16936 => "0000000000000000", 16937 => "0000000000000000", 16938 => "0000000000000000", 16939 => "0000000000000000", 16940 => "0000000000000000", 16941 => "0000000000000000", 16942 => "0000000000000000", 16943 => "0000000000000000", 16944 => "0000000000000000", 16945 => "0000000000000000", 16946 => "0000000000000000", 16947 => "0000000000000000", 16948 => "0000000000000000", 16949 => "0000000000000000", 16950 => "0000000000000000", 16951 => "0000000000000000", 16952 => "0000000000000000", 16953 => "0000000000000000", 16954 => "0000000000000000", 16955 => "0000000000000000", 16956 => "0000000000000000", 16957 => "0000000000000000", 16958 => "0000000000000000", 16959 => "0000000000000000", 16960 => "0000000000000000", 16961 => "0000000000000000", 16962 => "0000000000000000", 16963 => "0000000000000000", 16964 => "0000000000000000", 16965 => "0000000000000000", 16966 => "0000000000000000", 16967 => "0000000000000000", 16968 => "0000000000000000", 16969 => "0000000000000000", 16970 => "0000000000000000", 16971 => "0000000000000000", 16972 => "0000000000000000", 16973 => "0000000000000000", 16974 => "0000000000000000", 16975 => "0000000000000000", 16976 => "0000000000000000", 16977 => "0000000000000000", 16978 => "0000000000000000", 16979 => "0000000000000000", 16980 => "0000000000000000", 16981 => "0000000000000000", 16982 => "0000000000000000", 16983 => "0000000000000000", 16984 => "0000000000000000", 16985 => "0000000000000000", 16986 => "0000000000000000", 16987 => "0000000000000000", 16988 => "0000000000000000", 16989 => "0000000000000000", 16990 => "0000000000000000", 16991 => "0000000000000000", 16992 => "0000000000000000", 16993 => "0000000000000000", 16994 => "0000000000000000", 16995 => "0000000000000000", 16996 => "0000000000000000", 16997 => "0000000000000000", 16998 => "0000000000000000", 16999 => "0000000000000000", 17000 => "0000000000000000", 17001 => "0000000000000000", 17002 => "0000000000000000", 17003 => "0000000000000000", 17004 => "0000000000000000", 17005 => "0000000000000000", 17006 => "0000000000000000", 17007 => "0000000000000000", 17008 => "0000000000000000", 17009 => "0000000000000000", 17010 => "0000000000000000", 17011 => "0000000000000000", 17012 => "0000000000000000", 17013 => "0000000000000000", 17014 => "0000000000000000", 17015 => "0000000000000000", 17016 => "0000000000000000", 17017 => "0000000000000000", 17018 => "0000000000000000", 17019 => "0000000000000000", 17020 => "0000000000000000", 17021 => "0000000000000000", 17022 => "0000000000000000", 17023 => "0000000000000000", 17024 => "0000000000000000", 17025 => "0000000000000000", 17026 => "0000000000000000", 17027 => "0000000000000000", 17028 => "0000000000000000", 17029 => "0000000000000000", 17030 => "0000000000000000", 17031 => "0000000000000000", 17032 => "0000000000000000", 17033 => "0000000000000000", 17034 => "0000000000000000", 17035 => "0000000000000000", 17036 => "0000000000000000", 17037 => "0000000000000000", 17038 => "0000000000000000", 17039 => "0000000000000000", 17040 => "0000000000000000", 17041 => "0000000000000000", 17042 => "0000000000000000", 17043 => "0000000000000000", 17044 => "0000000000000000", 17045 => "0000000000000000", 17046 => "0000000000000000", 17047 => "0000000000000000", 17048 => "0000000000000000", 17049 => "0000000000000000", 17050 => "0000000000000000", 17051 => "0000000000000000", 17052 => "0000000000000000", 17053 => "0000000000000000", 17054 => "0000000000000000", 17055 => "0000000000000000", 17056 => "0000000000000000", 17057 => "0000000000000000", 17058 => "0000000000000000", 17059 => "0000000000000000", 17060 => "0000000000000000", 17061 => "0000000000000000", 17062 => "0000000000000000", 17063 => "0000000000000000", 17064 => "0000000000000000", 17065 => "0000000000000000", 17066 => "0000000000000000", 17067 => "0000000000000000", 17068 => "0000000000000000", 17069 => "0000000000000000", 17070 => "0000000000000000", 17071 => "0000000000000000", 17072 => "0000000000000000", 17073 => "0000000000000000", 17074 => "0000000000000000", 17075 => "0000000000000000", 17076 => "0000000000000000", 17077 => "0000000000000000", 17078 => "0000000000000000", 17079 => "0000000000000000", 17080 => "0000000000000000", 17081 => "0000000000000000", 17082 => "0000000000000000", 17083 => "0000000000000000", 17084 => "0000000000000000", 17085 => "0000000000000000", 17086 => "0000000000000000", 17087 => "0000000000000000", 17088 => "0000000000000000", 17089 => "0000000000000000", 17090 => "0000000000000000", 17091 => "0000000000000000", 17092 => "0000000000000000", 17093 => "0000000000000000", 17094 => "0000000000000000", 17095 => "0000000000000000", 17096 => "0000000000000000", 17097 => "0000000000000000", 17098 => "0000000000000000", 17099 => "0000000000000000", 17100 => "0000000000000000", 17101 => "0000000000000000", 17102 => "0000000000000000", 17103 => "0000000000000000", 17104 => "0000000000000000", 17105 => "0000000000000000", 17106 => "0000000000000000", 17107 => "0000000000000000", 17108 => "0000000000000000", 17109 => "0000000000000000", 17110 => "0000000000000000", 17111 => "0000000000000000", 17112 => "0000000000000000", 17113 => "0000000000000000", 17114 => "0000000000000000", 17115 => "0000000000000000", 17116 => "0000000000000000", 17117 => "0000000000000000", 17118 => "0000000000000000", 17119 => "0000000000000000", 17120 => "0000000000000000", 17121 => "0000000000000000", 17122 => "0000000000000000", 17123 => "0000000000000000", 17124 => "0000000000000000", 17125 => "0000000000000000", 17126 => "0000000000000000", 17127 => "0000000000000000", 17128 => "0000000000000000", 17129 => "0000000000000000", 17130 => "0000000000000000", 17131 => "0000000000000000", 17132 => "0000000000000000", 17133 => "0000000000000000", 17134 => "0000000000000000", 17135 => "0000000000000000", 17136 => "0000000000000000", 17137 => "0000000000000000", 17138 => "0000000000000000", 17139 => "0000000000000000", 17140 => "0000000000000000", 17141 => "0000000000000000", 17142 => "0000000000000000", 17143 => "0000000000000000", 17144 => "0000000000000000", 17145 => "0000000000000000", 17146 => "0000000000000000", 17147 => "0000000000000000", 17148 => "0000000000000000", 17149 => "0000000000000000", 17150 => "0000000000000000", 17151 => "0000000000000000", 17152 => "0000000000000000", 17153 => "0000000000000000", 17154 => "0000000000000000", 17155 => "0000000000000000", 17156 => "0000000000000000", 17157 => "0000000000000000", 17158 => "0000000000000000", 17159 => "0000000000000000", 17160 => "0000000000000000", 17161 => "0000000000000000", 17162 => "0000000000000000", 17163 => "0000000000000000", 17164 => "0000000000000000", 17165 => "0000000000000000", 17166 => "0000000000000000", 17167 => "0000000000000000", 17168 => "0000000000000000", 17169 => "0000000000000000", 17170 => "0000000000000000", 17171 => "0000000000000000", 17172 => "0000000000000000", 17173 => "0000000000000000", 17174 => "0000000000000000", 17175 => "0000000000000000", 17176 => "0000000000000000", 17177 => "0000000000000000", 17178 => "0000000000000000", 17179 => "0000000000000000", 17180 => "0000000000000000", 17181 => "0000000000000000", 17182 => "0000000000000000", 17183 => "0000000000000000", 17184 => "0000000000000000", 17185 => "0000000000000000", 17186 => "0000000000000000", 17187 => "0000000000000000", 17188 => "0000000000000000", 17189 => "0000000000000000", 17190 => "0000000000000000", 17191 => "0000000000000000", 17192 => "0000000000000000", 17193 => "0000000000000000", 17194 => "0000000000000000", 17195 => "0000000000000000", 17196 => "0000000000000000", 17197 => "0000000000000000", 17198 => "0000000000000000", 17199 => "0000000000000000", 17200 => "0000000000000000", 17201 => "0000000000000000", 17202 => "0000000000000000", 17203 => "0000000000000000", 17204 => "0000000000000000", 17205 => "0000000000000000", 17206 => "0000000000000000", 17207 => "0000000000000000", 17208 => "0000000000000000", 17209 => "0000000000000000", 17210 => "0000000000000000", 17211 => "0000000000000000", 17212 => "0000000000000000", 17213 => "0000000000000000", 17214 => "0000000000000000", 17215 => "0000000000000000", 17216 => "0000000000000000", 17217 => "0000000000000000", 17218 => "0000000000000000", 17219 => "0000000000000000", 17220 => "0000000000000000", 17221 => "0000000000000000", 17222 => "0000000000000000", 17223 => "0000000000000000", 17224 => "0000000000000000", 17225 => "0000000000000000", 17226 => "0000000000000000", 17227 => "0000000000000000", 17228 => "0000000000000000", 17229 => "0000000000000000", 17230 => "0000000000000000", 17231 => "0000000000000000", 17232 => "0000000000000000", 17233 => "0000000000000000", 17234 => "0000000000000000", 17235 => "0000000000000000", 17236 => "0000000000000000", 17237 => "0000000000000000", 17238 => "0000000000000000", 17239 => "0000000000000000", 17240 => "0000000000000000", 17241 => "0000000000000000", 17242 => "0000000000000000", 17243 => "0000000000000000", 17244 => "0000000000000000", 17245 => "0000000000000000", 17246 => "0000000000000000", 17247 => "0000000000000000", 17248 => "0000000000000000", 17249 => "0000000000000000", 17250 => "0000000000000000", 17251 => "0000000000000000", 17252 => "0000000000000000", 17253 => "0000000000000000", 17254 => "0000000000000000", 17255 => "0000000000000000", 17256 => "0000000000000000", 17257 => "0000000000000000", 17258 => "0000000000000000", 17259 => "0000000000000000", 17260 => "0000000000000000", 17261 => "0000000000000000", 17262 => "0000000000000000", 17263 => "0000000000000000", 17264 => "0000000000000000", 17265 => "0000000000000000", 17266 => "0000000000000000", 17267 => "0000000000000000", 17268 => "0000000000000000", 17269 => "0000000000000000", 17270 => "0000000000000000", 17271 => "0000000000000000", 17272 => "0000000000000000", 17273 => "0000000000000000", 17274 => "0000000000000000", 17275 => "0000000000000000", 17276 => "0000000000000000", 17277 => "0000000000000000", 17278 => "0000000000000000", 17279 => "0000000000000000", 17280 => "0000000000000000", 17281 => "0000000000000000", 17282 => "0000000000000000", 17283 => "0000000000000000", 17284 => "0000000000000000", 17285 => "0000000000000000", 17286 => "0000000000000000", 17287 => "0000000000000000", 17288 => "0000000000000000", 17289 => "0000000000000000", 17290 => "0000000000000000", 17291 => "0000000000000000", 17292 => "0000000000000000", 17293 => "0000000000000000", 17294 => "0000000000000000", 17295 => "0000000000000000", 17296 => "0000000000000000", 17297 => "0000000000000000", 17298 => "0000000000000000", 17299 => "0000000000000000", 17300 => "0000000000000000", 17301 => "0000000000000000", 17302 => "0000000000000000", 17303 => "0000000000000000", 17304 => "0000000000000000", 17305 => "0000000000000000", 17306 => "0000000000000000", 17307 => "0000000000000000", 17308 => "0000000000000000", 17309 => "0000000000000000", 17310 => "0000000000000000", 17311 => "0000000000000000", 17312 => "0000000000000000", 17313 => "0000000000000000", 17314 => "0000000000000000", 17315 => "0000000000000000", 17316 => "0000000000000000", 17317 => "0000000000000000", 17318 => "0000000000000000", 17319 => "0000000000000000", 17320 => "0000000000000000", 17321 => "0000000000000000", 17322 => "0000000000000000", 17323 => "0000000000000000", 17324 => "0000000000000000", 17325 => "0000000000000000", 17326 => "0000000000000000", 17327 => "0000000000000000", 17328 => "0000000000000000", 17329 => "0000000000000000", 17330 => "0000000000000000", 17331 => "0000000000000000", 17332 => "0000000000000000", 17333 => "0000000000000000", 17334 => "0000000000000000", 17335 => "0000000000000000", 17336 => "0000000000000000", 17337 => "0000000000000000", 17338 => "0000000000000000", 17339 => "0000000000000000", 17340 => "0000000000000000", 17341 => "0000000000000000", 17342 => "0000000000000000", 17343 => "0000000000000000", 17344 => "0000000000000000", 17345 => "0000000000000000", 17346 => "0000000000000000", 17347 => "0000000000000000", 17348 => "0000000000000000", 17349 => "0000000000000000", 17350 => "0000000000000000", 17351 => "0000000000000000", 17352 => "0000000000000000", 17353 => "0000000000000000", 17354 => "0000000000000000", 17355 => "0000000000000000", 17356 => "0000000000000000", 17357 => "0000000000000000", 17358 => "0000000000000000", 17359 => "0000000000000000", 17360 => "0000000000000000", 17361 => "0000000000000000", 17362 => "0000000000000000", 17363 => "0000000000000000", 17364 => "0000000000000000", 17365 => "0000000000000000", 17366 => "0000000000000000", 17367 => "0000000000000000", 17368 => "0000000000000000", 17369 => "0000000000000000", 17370 => "0000000000000000", 17371 => "0000000000000000", 17372 => "0000000000000000", 17373 => "0000000000000000", 17374 => "0000000000000000", 17375 => "0000000000000000", 17376 => "0000000000000000", 17377 => "0000000000000000", 17378 => "0000000000000000", 17379 => "0000000000000000", 17380 => "0000000000000000", 17381 => "0000000000000000", 17382 => "0000000000000000", 17383 => "0000000000000000", 17384 => "0000000000000000", 17385 => "0000000000000000", 17386 => "0000000000000000", 17387 => "0000000000000000", 17388 => "0000000000000000", 17389 => "0000000000000000", 17390 => "0000000000000000", 17391 => "0000000000000000", 17392 => "0000000000000000", 17393 => "0000000000000000", 17394 => "0000000000000000", 17395 => "0000000000000000", 17396 => "0000000000000000", 17397 => "0000000000000000", 17398 => "0000000000000000", 17399 => "0000000000000000", 17400 => "0000000000000000", 17401 => "0000000000000000", 17402 => "0000000000000000", 17403 => "0000000000000000", 17404 => "0000000000000000", 17405 => "0000000000000000", 17406 => "0000000000000000", 17407 => "0000000000000000", 17408 => "0000000000000000", 17409 => "0000000000000000", 17410 => "0000000000000000", 17411 => "0000000000000000", 17412 => "0000000000000000", 17413 => "0000000000000000", 17414 => "0000000000000000", 17415 => "0000000000000000", 17416 => "0000000000000000", 17417 => "0000000000000000", 17418 => "0000000000000000", 17419 => "0000000000000000", 17420 => "0000000000000000", 17421 => "0000000000000000", 17422 => "0000000000000000", 17423 => "0000000000000000", 17424 => "0000000000000000", 17425 => "0000000000000000", 17426 => "0000000000000000", 17427 => "0000000000000000", 17428 => "0000000000000000", 17429 => "0000000000000000", 17430 => "0000000000000000", 17431 => "0000000000000000", 17432 => "0000000000000000", 17433 => "0000000000000000", 17434 => "0000000000000000", 17435 => "0000000000000000", 17436 => "0000000000000000", 17437 => "0000000000000000", 17438 => "0000000000000000", 17439 => "0000000000000000", 17440 => "0000000000000000", 17441 => "0000000000000000", 17442 => "0000000000000000", 17443 => "0000000000000000", 17444 => "0000000000000000", 17445 => "0000000000000000", 17446 => "0000000000000000", 17447 => "0000000000000000", 17448 => "0000000000000000", 17449 => "0000000000000000", 17450 => "0000000000000000", 17451 => "0000000000000000", 17452 => "0000000000000000", 17453 => "0000000000000000", 17454 => "0000000000000000", 17455 => "0000000000000000", 17456 => "0000000000000000", 17457 => "0000000000000000", 17458 => "0000000000000000", 17459 => "0000000000000000", 17460 => "0000000000000000", 17461 => "0000000000000000", 17462 => "0000000000000000", 17463 => "0000000000000000", 17464 => "0000000000000000", 17465 => "0000000000000000", 17466 => "0000000000000000", 17467 => "0000000000000000", 17468 => "0000000000000000", 17469 => "0000000000000000", 17470 => "0000000000000000", 17471 => "0000000000000000", 17472 => "0000000000000000", 17473 => "0000000000000000", 17474 => "0000000000000000", 17475 => "0000000000000000", 17476 => "0000000000000000", 17477 => "0000000000000000", 17478 => "0000000000000000", 17479 => "0000000000000000", 17480 => "0000000000000000", 17481 => "0000000000000000", 17482 => "0000000000000000", 17483 => "0000000000000000", 17484 => "0000000000000000", 17485 => "0000000000000000", 17486 => "0000000000000000", 17487 => "0000000000000000", 17488 => "0000000000000000", 17489 => "0000000000000000", 17490 => "0000000000000000", 17491 => "0000000000000000", 17492 => "0000000000000000", 17493 => "0000000000000000", 17494 => "0000000000000000", 17495 => "0000000000000000", 17496 => "0000000000000000", 17497 => "0000000000000000", 17498 => "0000000000000000", 17499 => "0000000000000000", 17500 => "0000000000000000", 17501 => "0000000000000000", 17502 => "0000000000000000", 17503 => "0000000000000000", 17504 => "0000000000000000", 17505 => "0000000000000000", 17506 => "0000000000000000", 17507 => "0000000000000000", 17508 => "0000000000000000", 17509 => "0000000000000000", 17510 => "0000000000000000", 17511 => "0000000000000000", 17512 => "0000000000000000", 17513 => "0000000000000000", 17514 => "0000000000000000", 17515 => "0000000000000000", 17516 => "0000000000000000", 17517 => "0000000000000000", 17518 => "0000000000000000", 17519 => "0000000000000000", 17520 => "0000000000000000", 17521 => "0000000000000000", 17522 => "0000000000000000", 17523 => "0000000000000000", 17524 => "0000000000000000", 17525 => "0000000000000000", 17526 => "0000000000000000", 17527 => "0000000000000000", 17528 => "0000000000000000", 17529 => "0000000000000000", 17530 => "0000000000000000", 17531 => "0000000000000000", 17532 => "0000000000000000", 17533 => "0000000000000000", 17534 => "0000000000000000", 17535 => "0000000000000000", 17536 => "0000000000000000", 17537 => "0000000000000000", 17538 => "0000000000000000", 17539 => "0000000000000000", 17540 => "0000000000000000", 17541 => "0000000000000000", 17542 => "0000000000000000", 17543 => "0000000000000000", 17544 => "0000000000000000", 17545 => "0000000000000000", 17546 => "0000000000000000", 17547 => "0000000000000000", 17548 => "0000000000000000", 17549 => "0000000000000000", 17550 => "0000000000000000", 17551 => "0000000000000000", 17552 => "0000000000000000", 17553 => "0000000000000000", 17554 => "0000000000000000", 17555 => "0000000000000000", 17556 => "0000000000000000", 17557 => "0000000000000000", 17558 => "0000000000000000", 17559 => "0000000000000000", 17560 => "0000000000000000", 17561 => "0000000000000000", 17562 => "0000000000000000", 17563 => "0000000000000000", 17564 => "0000000000000000", 17565 => "0000000000000000", 17566 => "0000000000000000", 17567 => "0000000000000000", 17568 => "0000000000000000", 17569 => "0000000000000000", 17570 => "0000000000000000", 17571 => "0000000000000000", 17572 => "0000000000000000", 17573 => "0000000000000000", 17574 => "0000000000000000", 17575 => "0000000000000000", 17576 => "0000000000000000", 17577 => "0000000000000000", 17578 => "0000000000000000", 17579 => "0000000000000000", 17580 => "0000000000000000", 17581 => "0000000000000000", 17582 => "0000000000000000", 17583 => "0000000000000000", 17584 => "0000000000000000", 17585 => "0000000000000000", 17586 => "0000000000000000", 17587 => "0000000000000000", 17588 => "0000000000000000", 17589 => "0000000000000000", 17590 => "0000000000000000", 17591 => "0000000000000000", 17592 => "0000000000000000", 17593 => "0000000000000000", 17594 => "0000000000000000", 17595 => "0000000000000000", 17596 => "0000000000000000", 17597 => "0000000000000000", 17598 => "0000000000000000", 17599 => "0000000000000000", 17600 => "0000000000000000", 17601 => "0000000000000000", 17602 => "0000000000000000", 17603 => "0000000000000000", 17604 => "0000000000000000", 17605 => "0000000000000000", 17606 => "0000000000000000", 17607 => "0000000000000000", 17608 => "0000000000000000", 17609 => "0000000000000000", 17610 => "0000000000000000", 17611 => "0000000000000000", 17612 => "0000000000000000", 17613 => "0000000000000000", 17614 => "0000000000000000", 17615 => "0000000000000000", 17616 => "0000000000000000", 17617 => "0000000000000000", 17618 => "0000000000000000", 17619 => "0000000000000000", 17620 => "0000000000000000", 17621 => "0000000000000000", 17622 => "0000000000000000", 17623 => "0000000000000000", 17624 => "0000000000000000", 17625 => "0000000000000000", 17626 => "0000000000000000", 17627 => "0000000000000000", 17628 => "0000000000000000", 17629 => "0000000000000000", 17630 => "0000000000000000", 17631 => "0000000000000000", 17632 => "0000000000000000", 17633 => "0000000000000000", 17634 => "0000000000000000", 17635 => "0000000000000000", 17636 => "0000000000000000", 17637 => "0000000000000000", 17638 => "0000000000000000", 17639 => "0000000000000000", 17640 => "0000000000000000", 17641 => "0000000000000000", 17642 => "0000000000000000", 17643 => "0000000000000000", 17644 => "0000000000000000", 17645 => "0000000000000000", 17646 => "0000000000000000", 17647 => "0000000000000000", 17648 => "0000000000000000", 17649 => "0000000000000000", 17650 => "0000000000000000", 17651 => "0000000000000000", 17652 => "0000000000000000", 17653 => "0000000000000000", 17654 => "0000000000000000", 17655 => "0000000000000000", 17656 => "0000000000000000", 17657 => "0000000000000000", 17658 => "0000000000000000", 17659 => "0000000000000000", 17660 => "0000000000000000", 17661 => "0000000000000000", 17662 => "0000000000000000", 17663 => "0000000000000000", 17664 => "0000000000000000", 17665 => "0000000000000000", 17666 => "0000000000000000", 17667 => "0000000000000000", 17668 => "0000000000000000", 17669 => "0000000000000000", 17670 => "0000000000000000", 17671 => "0000000000000000", 17672 => "0000000000000000", 17673 => "0000000000000000", 17674 => "0000000000000000", 17675 => "0000000000000000", 17676 => "0000000000000000", 17677 => "0000000000000000", 17678 => "0000000000000000", 17679 => "0000000000000000", 17680 => "0000000000000000", 17681 => "0000000000000000", 17682 => "0000000000000000", 17683 => "0000000000000000", 17684 => "0000000000000000", 17685 => "0000000000000000", 17686 => "0000000000000000", 17687 => "0000000000000000", 17688 => "0000000000000000", 17689 => "0000000000000000", 17690 => "0000000000000000", 17691 => "0000000000000000", 17692 => "0000000000000000", 17693 => "0000000000000000", 17694 => "0000000000000000", 17695 => "0000000000000000", 17696 => "0000000000000000", 17697 => "0000000000000000", 17698 => "0000000000000000", 17699 => "0000000000000000", 17700 => "0000000000000000", 17701 => "0000000000000000", 17702 => "0000000000000000", 17703 => "0000000000000000", 17704 => "0000000000000000", 17705 => "0000000000000000", 17706 => "0000000000000000", 17707 => "0000000000000000", 17708 => "0000000000000000", 17709 => "0000000000000000", 17710 => "0000000000000000", 17711 => "0000000000000000", 17712 => "0000000000000000", 17713 => "0000000000000000", 17714 => "0000000000000000", 17715 => "0000000000000000", 17716 => "0000000000000000", 17717 => "0000000000000000", 17718 => "0000000000000000", 17719 => "0000000000000000", 17720 => "0000000000000000", 17721 => "0000000000000000", 17722 => "0000000000000000", 17723 => "0000000000000000", 17724 => "0000000000000000", 17725 => "0000000000000000", 17726 => "0000000000000000", 17727 => "0000000000000000", 17728 => "0000000000000000", 17729 => "0000000000000000", 17730 => "0000000000000000", 17731 => "0000000000000000", 17732 => "0000000000000000", 17733 => "0000000000000000", 17734 => "0000000000000000", 17735 => "0000000000000000", 17736 => "0000000000000000", 17737 => "0000000000000000", 17738 => "0000000000000000", 17739 => "0000000000000000", 17740 => "0000000000000000", 17741 => "0000000000000000", 17742 => "0000000000000000", 17743 => "0000000000000000", 17744 => "0000000000000000", 17745 => "0000000000000000", 17746 => "0000000000000000", 17747 => "0000000000000000", 17748 => "0000000000000000", 17749 => "0000000000000000", 17750 => "0000000000000000", 17751 => "0000000000000000", 17752 => "0000000000000000", 17753 => "0000000000000000", 17754 => "0000000000000000", 17755 => "0000000000000000", 17756 => "0000000000000000", 17757 => "0000000000000000", 17758 => "0000000000000000", 17759 => "0000000000000000", 17760 => "0000000000000000", 17761 => "0000000000000000", 17762 => "0000000000000000", 17763 => "0000000000000000", 17764 => "0000000000000000", 17765 => "0000000000000000", 17766 => "0000000000000000", 17767 => "0000000000000000", 17768 => "0000000000000000", 17769 => "0000000000000000", 17770 => "0000000000000000", 17771 => "0000000000000000", 17772 => "0000000000000000", 17773 => "0000000000000000", 17774 => "0000000000000000", 17775 => "0000000000000000", 17776 => "0000000000000000", 17777 => "0000000000000000", 17778 => "0000000000000000", 17779 => "0000000000000000", 17780 => "0000000000000000", 17781 => "0000000000000000", 17782 => "0000000000000000", 17783 => "0000000000000000", 17784 => "0000000000000000", 17785 => "0000000000000000", 17786 => "0000000000000000", 17787 => "0000000000000000", 17788 => "0000000000000000", 17789 => "0000000000000000", 17790 => "0000000000000000", 17791 => "0000000000000000", 17792 => "0000000000000000", 17793 => "0000000000000000", 17794 => "0000000000000000", 17795 => "0000000000000000", 17796 => "0000000000000000", 17797 => "0000000000000000", 17798 => "0000000000000000", 17799 => "0000000000000000", 17800 => "0000000000000000", 17801 => "0000000000000000", 17802 => "0000000000000000", 17803 => "0000000000000000", 17804 => "0000000000000000", 17805 => "0000000000000000", 17806 => "0000000000000000", 17807 => "0000000000000000", 17808 => "0000000000000000", 17809 => "0000000000000000", 17810 => "0000000000000000", 17811 => "0000000000000000", 17812 => "0000000000000000", 17813 => "0000000000000000", 17814 => "0000000000000000", 17815 => "0000000000000000", 17816 => "0000000000000000", 17817 => "0000000000000000", 17818 => "0000000000000000", 17819 => "0000000000000000", 17820 => "0000000000000000", 17821 => "0000000000000000", 17822 => "0000000000000000", 17823 => "0000000000000000", 17824 => "0000000000000000", 17825 => "0000000000000000", 17826 => "0000000000000000", 17827 => "0000000000000000", 17828 => "0000000000000000", 17829 => "0000000000000000", 17830 => "0000000000000000", 17831 => "0000000000000000", 17832 => "0000000000000000", 17833 => "0000000000000000", 17834 => "0000000000000000", 17835 => "0000000000000000", 17836 => "0000000000000000", 17837 => "0000000000000000", 17838 => "0000000000000000", 17839 => "0000000000000000", 17840 => "0000000000000000", 17841 => "0000000000000000", 17842 => "0000000000000000", 17843 => "0000000000000000", 17844 => "0000000000000000", 17845 => "0000000000000000", 17846 => "0000000000000000", 17847 => "0000000000000000", 17848 => "0000000000000000", 17849 => "0000000000000000", 17850 => "0000000000000000", 17851 => "0000000000000000", 17852 => "0000000000000000", 17853 => "0000000000000000", 17854 => "0000000000000000", 17855 => "0000000000000000", 17856 => "0000000000000000", 17857 => "0000000000000000", 17858 => "0000000000000000", 17859 => "0000000000000000", 17860 => "0000000000000000", 17861 => "0000000000000000", 17862 => "0000000000000000", 17863 => "0000000000000000", 17864 => "0000000000000000", 17865 => "0000000000000000", 17866 => "0000000000000000", 17867 => "0000000000000000", 17868 => "0000000000000000", 17869 => "0000000000000000", 17870 => "0000000000000000", 17871 => "0000000000000000", 17872 => "0000000000000000", 17873 => "0000000000000000", 17874 => "0000000000000000", 17875 => "0000000000000000", 17876 => "0000000000000000", 17877 => "0000000000000000", 17878 => "0000000000000000", 17879 => "0000000000000000", 17880 => "0000000000000000", 17881 => "0000000000000000", 17882 => "0000000000000000", 17883 => "0000000000000000", 17884 => "0000000000000000", 17885 => "0000000000000000", 17886 => "0000000000000000", 17887 => "0000000000000000", 17888 => "0000000000000000", 17889 => "0000000000000000", 17890 => "0000000000000000", 17891 => "0000000000000000", 17892 => "0000000000000000", 17893 => "0000000000000000", 17894 => "0000000000000000", 17895 => "0000000000000000", 17896 => "0000000000000000", 17897 => "0000000000000000", 17898 => "0000000000000000", 17899 => "0000000000000000", 17900 => "0000000000000000", 17901 => "0000000000000000", 17902 => "0000000000000000", 17903 => "0000000000000000", 17904 => "0000000000000000", 17905 => "0000000000000000", 17906 => "0000000000000000", 17907 => "0000000000000000", 17908 => "0000000000000000", 17909 => "0000000000000000", 17910 => "0000000000000000", 17911 => "0000000000000000", 17912 => "0000000000000000", 17913 => "0000000000000000", 17914 => "0000000000000000", 17915 => "0000000000000000", 17916 => "0000000000000000", 17917 => "0000000000000000", 17918 => "0000000000000000", 17919 => "0000000000000000", 17920 => "0000000000000000", 17921 => "0000000000000000", 17922 => "0000000000000000", 17923 => "0000000000000000", 17924 => "0000000000000000", 17925 => "0000000000000000", 17926 => "0000000000000000", 17927 => "0000000000000000", 17928 => "0000000000000000", 17929 => "0000000000000000", 17930 => "0000000000000000", 17931 => "0000000000000000", 17932 => "0000000000000000", 17933 => "0000000000000000", 17934 => "0000000000000000", 17935 => "0000000000000000", 17936 => "0000000000000000", 17937 => "0000000000000000", 17938 => "0000000000000000", 17939 => "0000000000000000", 17940 => "0000000000000000", 17941 => "0000000000000000", 17942 => "0000000000000000", 17943 => "0000000000000000", 17944 => "0000000000000000", 17945 => "0000000000000000", 17946 => "0000000000000000", 17947 => "0000000000000000", 17948 => "0000000000000000", 17949 => "0000000000000000", 17950 => "0000000000000000", 17951 => "0000000000000000", 17952 => "0000000000000000", 17953 => "0000000000000000", 17954 => "0000000000000000", 17955 => "0000000000000000", 17956 => "0000000000000000", 17957 => "0000000000000000", 17958 => "0000000000000000", 17959 => "0000000000000000", 17960 => "0000000000000000", 17961 => "0000000000000000", 17962 => "0000000000000000", 17963 => "0000000000000000", 17964 => "0000000000000000", 17965 => "0000000000000000", 17966 => "0000000000000000", 17967 => "0000000000000000", 17968 => "0000000000000000", 17969 => "0000000000000000", 17970 => "0000000000000000", 17971 => "0000000000000000", 17972 => "0000000000000000", 17973 => "0000000000000000", 17974 => "0000000000000000", 17975 => "0000000000000000", 17976 => "0000000000000000", 17977 => "0000000000000000", 17978 => "0000000000000000", 17979 => "0000000000000000", 17980 => "0000000000000000", 17981 => "0000000000000000", 17982 => "0000000000000000", 17983 => "0000000000000000", 17984 => "0000000000000000", 17985 => "0000000000000000", 17986 => "0000000000000000", 17987 => "0000000000000000", 17988 => "0000000000000000", 17989 => "0000000000000000", 17990 => "0000000000000000", 17991 => "0000000000000000", 17992 => "0000000000000000", 17993 => "0000000000000000", 17994 => "0000000000000000", 17995 => "0000000000000000", 17996 => "0000000000000000", 17997 => "0000000000000000", 17998 => "0000000000000000", 17999 => "0000000000000000", 18000 => "0000000000000000", 18001 => "0000000000000000", 18002 => "0000000000000000", 18003 => "0000000000000000", 18004 => "0000000000000000", 18005 => "0000000000000000", 18006 => "0000000000000000", 18007 => "0000000000000000", 18008 => "0000000000000000", 18009 => "0000000000000000", 18010 => "0000000000000000", 18011 => "0000000000000000", 18012 => "0000000000000000", 18013 => "0000000000000000", 18014 => "0000000000000000", 18015 => "0000000000000000", 18016 => "0000000000000000", 18017 => "0000000000000000", 18018 => "0000000000000000", 18019 => "0000000000000000", 18020 => "0000000000000000", 18021 => "0000000000000000", 18022 => "0000000000000000", 18023 => "0000000000000000", 18024 => "0000000000000000", 18025 => "0000000000000000", 18026 => "0000000000000000", 18027 => "0000000000000000", 18028 => "0000000000000000", 18029 => "0000000000000000", 18030 => "0000000000000000", 18031 => "0000000000000000", 18032 => "0000000000000000", 18033 => "0000000000000000", 18034 => "0000000000000000", 18035 => "0000000000000000", 18036 => "0000000000000000", 18037 => "0000000000000000", 18038 => "0000000000000000", 18039 => "0000000000000000", 18040 => "0000000000000000", 18041 => "0000000000000000", 18042 => "0000000000000000", 18043 => "0000000000000000", 18044 => "0000000000000000", 18045 => "0000000000000000", 18046 => "0000000000000000", 18047 => "0000000000000000", 18048 => "0000000000000000", 18049 => "0000000000000000", 18050 => "0000000000000000", 18051 => "0000000000000000", 18052 => "0000000000000000", 18053 => "0000000000000000", 18054 => "0000000000000000", 18055 => "0000000000000000", 18056 => "0000000000000000", 18057 => "0000000000000000", 18058 => "0000000000000000", 18059 => "0000000000000000", 18060 => "0000000000000000", 18061 => "0000000000000000", 18062 => "0000000000000000", 18063 => "0000000000000000", 18064 => "0000000000000000", 18065 => "0000000000000000", 18066 => "0000000000000000", 18067 => "0000000000000000", 18068 => "0000000000000000", 18069 => "0000000000000000", 18070 => "0000000000000000", 18071 => "0000000000000000", 18072 => "0000000000000000", 18073 => "0000000000000000", 18074 => "0000000000000000", 18075 => "0000000000000000", 18076 => "0000000000000000", 18077 => "0000000000000000", 18078 => "0000000000000000", 18079 => "0000000000000000", 18080 => "0000000000000000", 18081 => "0000000000000000", 18082 => "0000000000000000", 18083 => "0000000000000000", 18084 => "0000000000000000", 18085 => "0000000000000000", 18086 => "0000000000000000", 18087 => "0000000000000000", 18088 => "0000000000000000", 18089 => "0000000000000000", 18090 => "0000000000000000", 18091 => "0000000000000000", 18092 => "0000000000000000", 18093 => "0000000000000000", 18094 => "0000000000000000", 18095 => "0000000000000000", 18096 => "0000000000000000", 18097 => "0000000000000000", 18098 => "0000000000000000", 18099 => "0000000000000000", 18100 => "0000000000000000", 18101 => "0000000000000000", 18102 => "0000000000000000", 18103 => "0000000000000000", 18104 => "0000000000000000", 18105 => "0000000000000000", 18106 => "0000000000000000", 18107 => "0000000000000000", 18108 => "0000000000000000", 18109 => "0000000000000000", 18110 => "0000000000000000", 18111 => "0000000000000000", 18112 => "0000000000000000", 18113 => "0000000000000000", 18114 => "0000000000000000", 18115 => "0000000000000000", 18116 => "0000000000000000", 18117 => "0000000000000000", 18118 => "0000000000000000", 18119 => "0000000000000000", 18120 => "0000000000000000", 18121 => "0000000000000000", 18122 => "0000000000000000", 18123 => "0000000000000000", 18124 => "0000000000000000", 18125 => "0000000000000000", 18126 => "0000000000000000", 18127 => "0000000000000000", 18128 => "0000000000000000", 18129 => "0000000000000000", 18130 => "0000000000000000", 18131 => "0000000000000000", 18132 => "0000000000000000", 18133 => "0000000000000000", 18134 => "0000000000000000", 18135 => "0000000000000000", 18136 => "0000000000000000", 18137 => "0000000000000000", 18138 => "0000000000000000", 18139 => "0000000000000000", 18140 => "0000000000000000", 18141 => "0000000000000000", 18142 => "0000000000000000", 18143 => "0000000000000000", 18144 => "0000000000000000", 18145 => "0000000000000000", 18146 => "0000000000000000", 18147 => "0000000000000000", 18148 => "0000000000000000", 18149 => "0000000000000000", 18150 => "0000000000000000", 18151 => "0000000000000000", 18152 => "0000000000000000", 18153 => "0000000000000000", 18154 => "0000000000000000", 18155 => "0000000000000000", 18156 => "0000000000000000", 18157 => "0000000000000000", 18158 => "0000000000000000", 18159 => "0000000000000000", 18160 => "0000000000000000", 18161 => "0000000000000000", 18162 => "0000000000000000", 18163 => "0000000000000000", 18164 => "0000000000000000", 18165 => "0000000000000000", 18166 => "0000000000000000", 18167 => "0000000000000000", 18168 => "0000000000000000", 18169 => "0000000000000000", 18170 => "0000000000000000", 18171 => "0000000000000000", 18172 => "0000000000000000", 18173 => "0000000000000000", 18174 => "0000000000000000", 18175 => "0000000000000000", 18176 => "0000000000000000", 18177 => "0000000000000000", 18178 => "0000000000000000", 18179 => "0000000000000000", 18180 => "0000000000000000", 18181 => "0000000000000000", 18182 => "0000000000000000", 18183 => "0000000000000000", 18184 => "0000000000000000", 18185 => "0000000000000000", 18186 => "0000000000000000", 18187 => "0000000000000000", 18188 => "0000000000000000", 18189 => "0000000000000000", 18190 => "0000000000000000", 18191 => "0000000000000000", 18192 => "0000000000000000", 18193 => "0000000000000000", 18194 => "0000000000000000", 18195 => "0000000000000000", 18196 => "0000000000000000", 18197 => "0000000000000000", 18198 => "0000000000000000", 18199 => "0000000000000000", 18200 => "0000000000000000", 18201 => "0000000000000000", 18202 => "0000000000000000", 18203 => "0000000000000000", 18204 => "0000000000000000", 18205 => "0000000000000000", 18206 => "0000000000000000", 18207 => "0000000000000000", 18208 => "0000000000000000", 18209 => "0000000000000000", 18210 => "0000000000000000", 18211 => "0000000000000000", 18212 => "0000000000000000", 18213 => "0000000000000000", 18214 => "0000000000000000", 18215 => "0000000000000000", 18216 => "0000000000000000", 18217 => "0000000000000000", 18218 => "0000000000000000", 18219 => "0000000000000000", 18220 => "0000000000000000", 18221 => "0000000000000000", 18222 => "0000000000000000", 18223 => "0000000000000000", 18224 => "0000000000000000", 18225 => "0000000000000000", 18226 => "0000000000000000", 18227 => "0000000000000000", 18228 => "0000000000000000", 18229 => "0000000000000000", 18230 => "0000000000000000", 18231 => "0000000000000000", 18232 => "0000000000000000", 18233 => "0000000000000000", 18234 => "0000000000000000", 18235 => "0000000000000000", 18236 => "0000000000000000", 18237 => "0000000000000000", 18238 => "0000000000000000", 18239 => "0000000000000000", 18240 => "0000000000000000", 18241 => "0000000000000000", 18242 => "0000000000000000", 18243 => "0000000000000000", 18244 => "0000000000000000", 18245 => "0000000000000000", 18246 => "0000000000000000", 18247 => "0000000000000000", 18248 => "0000000000000000", 18249 => "0000000000000000", 18250 => "0000000000000000", 18251 => "0000000000000000", 18252 => "0000000000000000", 18253 => "0000000000000000", 18254 => "0000000000000000", 18255 => "0000000000000000", 18256 => "0000000000000000", 18257 => "0000000000000000", 18258 => "0000000000000000", 18259 => "0000000000000000", 18260 => "0000000000000000", 18261 => "0000000000000000", 18262 => "0000000000000000", 18263 => "0000000000000000", 18264 => "0000000000000000", 18265 => "0000000000000000", 18266 => "0000000000000000", 18267 => "0000000000000000", 18268 => "0000000000000000", 18269 => "0000000000000000", 18270 => "0000000000000000", 18271 => "0000000000000000", 18272 => "0000000000000000", 18273 => "0000000000000000", 18274 => "0000000000000000", 18275 => "0000000000000000", 18276 => "0000000000000000", 18277 => "0000000000000000", 18278 => "0000000000000000", 18279 => "0000000000000000", 18280 => "0000000000000000", 18281 => "0000000000000000", 18282 => "0000000000000000", 18283 => "0000000000000000", 18284 => "0000000000000000", 18285 => "0000000000000000", 18286 => "0000000000000000", 18287 => "0000000000000000", 18288 => "0000000000000000", 18289 => "0000000000000000", 18290 => "0000000000000000", 18291 => "0000000000000000", 18292 => "0000000000000000", 18293 => "0000000000000000", 18294 => "0000000000000000", 18295 => "0000000000000000", 18296 => "0000000000000000", 18297 => "0000000000000000", 18298 => "0000000000000000", 18299 => "0000000000000000", 18300 => "0000000000000000", 18301 => "0000000000000000", 18302 => "0000000000000000", 18303 => "0000000000000000", 18304 => "0000000000000000", 18305 => "0000000000000000", 18306 => "0000000000000000", 18307 => "0000000000000000", 18308 => "0000000000000000", 18309 => "0000000000000000", 18310 => "0000000000000000", 18311 => "0000000000000000", 18312 => "0000000000000000", 18313 => "0000000000000000", 18314 => "0000000000000000", 18315 => "0000000000000000", 18316 => "0000000000000000", 18317 => "0000000000000000", 18318 => "0000000000000000", 18319 => "0000000000000000", 18320 => "0000000000000000", 18321 => "0000000000000000", 18322 => "0000000000000000", 18323 => "0000000000000000", 18324 => "0000000000000000", 18325 => "0000000000000000", 18326 => "0000000000000000", 18327 => "0000000000000000", 18328 => "0000000000000000", 18329 => "0000000000000000", 18330 => "0000000000000000", 18331 => "0000000000000000", 18332 => "0000000000000000", 18333 => "0000000000000000", 18334 => "0000000000000000", 18335 => "0000000000000000", 18336 => "0000000000000000", 18337 => "0000000000000000", 18338 => "0000000000000000", 18339 => "0000000000000000", 18340 => "0000000000000000", 18341 => "0000000000000000", 18342 => "0000000000000000", 18343 => "0000000000000000", 18344 => "0000000000000000", 18345 => "0000000000000000", 18346 => "0000000000000000", 18347 => "0000000000000000", 18348 => "0000000000000000", 18349 => "0000000000000000", 18350 => "0000000000000000", 18351 => "0000000000000000", 18352 => "0000000000000000", 18353 => "0000000000000000", 18354 => "0000000000000000", 18355 => "0000000000000000", 18356 => "0000000000000000", 18357 => "0000000000000000", 18358 => "0000000000000000", 18359 => "0000000000000000", 18360 => "0000000000000000", 18361 => "0000000000000000", 18362 => "0000000000000000", 18363 => "0000000000000000", 18364 => "0000000000000000", 18365 => "0000000000000000", 18366 => "0000000000000000", 18367 => "0000000000000000", 18368 => "0000000000000000", 18369 => "0000000000000000", 18370 => "0000000000000000", 18371 => "0000000000000000", 18372 => "0000000000000000", 18373 => "0000000000000000", 18374 => "0000000000000000", 18375 => "0000000000000000", 18376 => "0000000000000000", 18377 => "0000000000000000", 18378 => "0000000000000000", 18379 => "0000000000000000", 18380 => "0000000000000000", 18381 => "0000000000000000", 18382 => "0000000000000000", 18383 => "0000000000000000", 18384 => "0000000000000000", 18385 => "0000000000000000", 18386 => "0000000000000000", 18387 => "0000000000000000", 18388 => "0000000000000000", 18389 => "0000000000000000", 18390 => "0000000000000000", 18391 => "0000000000000000", 18392 => "0000000000000000", 18393 => "0000000000000000", 18394 => "0000000000000000", 18395 => "0000000000000000", 18396 => "0000000000000000", 18397 => "0000000000000000", 18398 => "0000000000000000", 18399 => "0000000000000000", 18400 => "0000000000000000", 18401 => "0000000000000000", 18402 => "0000000000000000", 18403 => "0000000000000000", 18404 => "0000000000000000", 18405 => "0000000000000000", 18406 => "0000000000000000", 18407 => "0000000000000000", 18408 => "0000000000000000", 18409 => "0000000000000000", 18410 => "0000000000000000", 18411 => "0000000000000000", 18412 => "0000000000000000", 18413 => "0000000000000000", 18414 => "0000000000000000", 18415 => "0000000000000000", 18416 => "0000000000000000", 18417 => "0000000000000000", 18418 => "0000000000000000", 18419 => "0000000000000000", 18420 => "0000000000000000", 18421 => "0000000000000000", 18422 => "0000000000000000", 18423 => "0000000000000000", 18424 => "0000000000000000", 18425 => "0000000000000000", 18426 => "0000000000000000", 18427 => "0000000000000000", 18428 => "0000000000000000", 18429 => "0000000000000000", 18430 => "0000000000000000", 18431 => "0000000000000000", 18432 => "0000000000000000", 18433 => "0000000000000000", 18434 => "0000000000000000", 18435 => "0000000000000000", 18436 => "0000000000000000", 18437 => "0000000000000000", 18438 => "0000000000000000", 18439 => "0000000000000000", 18440 => "0000000000000000", 18441 => "0000000000000000", 18442 => "0000000000000000", 18443 => "0000000000000000", 18444 => "0000000000000000", 18445 => "0000000000000000", 18446 => "0000000000000000", 18447 => "0000000000000000", 18448 => "0000000000000000", 18449 => "0000000000000000", 18450 => "0000000000000000", 18451 => "0000000000000000", 18452 => "0000000000000000", 18453 => "0000000000000000", 18454 => "0000000000000000", 18455 => "0000000000000000", 18456 => "0000000000000000", 18457 => "0000000000000000", 18458 => "0000000000000000", 18459 => "0000000000000000", 18460 => "0000000000000000", 18461 => "0000000000000000", 18462 => "0000000000000000", 18463 => "0000000000000000", 18464 => "0000000000000000", 18465 => "0000000000000000", 18466 => "0000000000000000", 18467 => "0000000000000000", 18468 => "0000000000000000", 18469 => "0000000000000000", 18470 => "0000000000000000", 18471 => "0000000000000000", 18472 => "0000000000000000", 18473 => "0000000000000000", 18474 => "0000000000000000", 18475 => "0000000000000000", 18476 => "0000000000000000", 18477 => "0000000000000000", 18478 => "0000000000000000", 18479 => "0000000000000000", 18480 => "0000000000000000", 18481 => "0000000000000000", 18482 => "0000000000000000", 18483 => "0000000000000000", 18484 => "0000000000000000", 18485 => "0000000000000000", 18486 => "0000000000000000", 18487 => "0000000000000000", 18488 => "0000000000000000", 18489 => "0000000000000000", 18490 => "0000000000000000", 18491 => "0000000000000000", 18492 => "0000000000000000", 18493 => "0000000000000000", 18494 => "0000000000000000", 18495 => "0000000000000000", 18496 => "0000000000000000", 18497 => "0000000000000000", 18498 => "0000000000000000", 18499 => "0000000000000000", 18500 => "0000000000000000", 18501 => "0000000000000000", 18502 => "0000000000000000", 18503 => "0000000000000000", 18504 => "0000000000000000", 18505 => "0000000000000000", 18506 => "0000000000000000", 18507 => "0000000000000000", 18508 => "0000000000000000", 18509 => "0000000000000000", 18510 => "0000000000000000", 18511 => "0000000000000000", 18512 => "0000000000000000", 18513 => "0000000000000000", 18514 => "0000000000000000", 18515 => "0000000000000000", 18516 => "0000000000000000", 18517 => "0000000000000000", 18518 => "0000000000000000", 18519 => "0000000000000000", 18520 => "0000000000000000", 18521 => "0000000000000000", 18522 => "0000000000000000", 18523 => "0000000000000000", 18524 => "0000000000000000", 18525 => "0000000000000000", 18526 => "0000000000000000", 18527 => "0000000000000000", 18528 => "0000000000000000", 18529 => "0000000000000000", 18530 => "0000000000000000", 18531 => "0000000000000000", 18532 => "0000000000000000", 18533 => "0000000000000000", 18534 => "0000000000000000", 18535 => "0000000000000000", 18536 => "0000000000000000", 18537 => "0000000000000000", 18538 => "0000000000000000", 18539 => "0000000000000000", 18540 => "0000000000000000", 18541 => "0000000000000000", 18542 => "0000000000000000", 18543 => "0000000000000000", 18544 => "0000000000000000", 18545 => "0000000000000000", 18546 => "0000000000000000", 18547 => "0000000000000000", 18548 => "0000000000000000", 18549 => "0000000000000000", 18550 => "0000000000000000", 18551 => "0000000000000000", 18552 => "0000000000000000", 18553 => "0000000000000000", 18554 => "0000000000000000", 18555 => "0000000000000000", 18556 => "0000000000000000", 18557 => "0000000000000000", 18558 => "0000000000000000", 18559 => "0000000000000000", 18560 => "0000000000000000", 18561 => "0000000000000000", 18562 => "0000000000000000", 18563 => "0000000000000000", 18564 => "0000000000000000", 18565 => "0000000000000000", 18566 => "0000000000000000", 18567 => "0000000000000000", 18568 => "0000000000000000", 18569 => "0000000000000000", 18570 => "0000000000000000", 18571 => "0000000000000000", 18572 => "0000000000000000", 18573 => "0000000000000000", 18574 => "0000000000000000", 18575 => "0000000000000000", 18576 => "0000000000000000", 18577 => "0000000000000000", 18578 => "0000000000000000", 18579 => "0000000000000000", 18580 => "0000000000000000", 18581 => "0000000000000000", 18582 => "0000000000000000", 18583 => "0000000000000000", 18584 => "0000000000000000", 18585 => "0000000000000000", 18586 => "0000000000000000", 18587 => "0000000000000000", 18588 => "0000000000000000", 18589 => "0000000000000000", 18590 => "0000000000000000", 18591 => "0000000000000000", 18592 => "0000000000000000", 18593 => "0000000000000000", 18594 => "0000000000000000", 18595 => "0000000000000000", 18596 => "0000000000000000", 18597 => "0000000000000000", 18598 => "0000000000000000", 18599 => "0000000000000000", 18600 => "0000000000000000", 18601 => "0000000000000000", 18602 => "0000000000000000", 18603 => "0000000000000000", 18604 => "0000000000000000", 18605 => "0000000000000000", 18606 => "0000000000000000", 18607 => "0000000000000000", 18608 => "0000000000000000", 18609 => "0000000000000000", 18610 => "0000000000000000", 18611 => "0000000000000000", 18612 => "0000000000000000", 18613 => "0000000000000000", 18614 => "0000000000000000", 18615 => "0000000000000000", 18616 => "0000000000000000", 18617 => "0000000000000000", 18618 => "0000000000000000", 18619 => "0000000000000000", 18620 => "0000000000000000", 18621 => "0000000000000000", 18622 => "0000000000000000", 18623 => "0000000000000000", 18624 => "0000000000000000", 18625 => "0000000000000000", 18626 => "0000000000000000", 18627 => "0000000000000000", 18628 => "0000000000000000", 18629 => "0000000000000000", 18630 => "0000000000000000", 18631 => "0000000000000000", 18632 => "0000000000000000", 18633 => "0000000000000000", 18634 => "0000000000000000", 18635 => "0000000000000000", 18636 => "0000000000000000", 18637 => "0000000000000000", 18638 => "0000000000000000", 18639 => "0000000000000000", 18640 => "0000000000000000", 18641 => "0000000000000000", 18642 => "0000000000000000", 18643 => "0000000000000000", 18644 => "0000000000000000", 18645 => "0000000000000000", 18646 => "0000000000000000", 18647 => "0000000000000000", 18648 => "0000000000000000", 18649 => "0000000000000000", 18650 => "0000000000000000", 18651 => "0000000000000000", 18652 => "0000000000000000", 18653 => "0000000000000000", 18654 => "0000000000000000", 18655 => "0000000000000000", 18656 => "0000000000000000", 18657 => "0000000000000000", 18658 => "0000000000000000", 18659 => "0000000000000000", 18660 => "0000000000000000", 18661 => "0000000000000000", 18662 => "0000000000000000", 18663 => "0000000000000000", 18664 => "0000000000000000", 18665 => "0000000000000000", 18666 => "0000000000000000", 18667 => "0000000000000000", 18668 => "0000000000000000", 18669 => "0000000000000000", 18670 => "0000000000000000", 18671 => "0000000000000000", 18672 => "0000000000000000", 18673 => "0000000000000000", 18674 => "0000000000000000", 18675 => "0000000000000000", 18676 => "0000000000000000", 18677 => "0000000000000000", 18678 => "0000000000000000", 18679 => "0000000000000000", 18680 => "0000000000000000", 18681 => "0000000000000000", 18682 => "0000000000000000", 18683 => "0000000000000000", 18684 => "0000000000000000", 18685 => "0000000000000000", 18686 => "0000000000000000", 18687 => "0000000000000000", 18688 => "0000000000000000", 18689 => "0000000000000000", 18690 => "0000000000000000", 18691 => "0000000000000000", 18692 => "0000000000000000", 18693 => "0000000000000000", 18694 => "0000000000000000", 18695 => "0000000000000000", 18696 => "0000000000000000", 18697 => "0000000000000000", 18698 => "0000000000000000", 18699 => "0000000000000000", 18700 => "0000000000000000", 18701 => "0000000000000000", 18702 => "0000000000000000", 18703 => "0000000000000000", 18704 => "0000000000000000", 18705 => "0000000000000000", 18706 => "0000000000000000", 18707 => "0000000000000000", 18708 => "0000000000000000", 18709 => "0000000000000000", 18710 => "0000000000000000", 18711 => "0000000000000000", 18712 => "0000000000000000", 18713 => "0000000000000000", 18714 => "0000000000000000", 18715 => "0000000000000000", 18716 => "0000000000000000", 18717 => "0000000000000000", 18718 => "0000000000000000", 18719 => "0000000000000000", 18720 => "0000000000000000", 18721 => "0000000000000000", 18722 => "0000000000000000", 18723 => "0000000000000000", 18724 => "0000000000000000", 18725 => "0000000000000000", 18726 => "0000000000000000", 18727 => "0000000000000000", 18728 => "0000000000000000", 18729 => "0000000000000000", 18730 => "0000000000000000", 18731 => "0000000000000000", 18732 => "0000000000000000", 18733 => "0000000000000000", 18734 => "0000000000000000", 18735 => "0000000000000000", 18736 => "0000000000000000", 18737 => "0000000000000000", 18738 => "0000000000000000", 18739 => "0000000000000000", 18740 => "0000000000000000", 18741 => "0000000000000000", 18742 => "0000000000000000", 18743 => "0000000000000000", 18744 => "0000000000000000", 18745 => "0000000000000000", 18746 => "0000000000000000", 18747 => "0000000000000000", 18748 => "0000000000000000", 18749 => "0000000000000000", 18750 => "0000000000000000", 18751 => "0000000000000000", 18752 => "0000000000000000", 18753 => "0000000000000000", 18754 => "0000000000000000", 18755 => "0000000000000000", 18756 => "0000000000000000", 18757 => "0000000000000000", 18758 => "0000000000000000", 18759 => "0000000000000000", 18760 => "0000000000000000", 18761 => "0000000000000000", 18762 => "0000000000000000", 18763 => "0000000000000000", 18764 => "0000000000000000", 18765 => "0000000000000000", 18766 => "0000000000000000", 18767 => "0000000000000000", 18768 => "0000000000000000", 18769 => "0000000000000000", 18770 => "0000000000000000", 18771 => "0000000000000000", 18772 => "0000000000000000", 18773 => "0000000000000000", 18774 => "0000000000000000", 18775 => "0000000000000000", 18776 => "0000000000000000", 18777 => "0000000000000000", 18778 => "0000000000000000", 18779 => "0000000000000000", 18780 => "0000000000000000", 18781 => "0000000000000000", 18782 => "0000000000000000", 18783 => "0000000000000000", 18784 => "0000000000000000", 18785 => "0000000000000000", 18786 => "0000000000000000", 18787 => "0000000000000000", 18788 => "0000000000000000", 18789 => "0000000000000000", 18790 => "0000000000000000", 18791 => "0000000000000000", 18792 => "0000000000000000", 18793 => "0000000000000000", 18794 => "0000000000000000", 18795 => "0000000000000000", 18796 => "0000000000000000", 18797 => "0000000000000000", 18798 => "0000000000000000", 18799 => "0000000000000000", 18800 => "0000000000000000", 18801 => "0000000000000000", 18802 => "0000000000000000", 18803 => "0000000000000000", 18804 => "0000000000000000", 18805 => "0000000000000000", 18806 => "0000000000000000", 18807 => "0000000000000000", 18808 => "0000000000000000", 18809 => "0000000000000000", 18810 => "0000000000000000", 18811 => "0000000000000000", 18812 => "0000000000000000", 18813 => "0000000000000000", 18814 => "0000000000000000", 18815 => "0000000000000000", 18816 => "0000000000000000", 18817 => "0000000000000000", 18818 => "0000000000000000", 18819 => "0000000000000000", 18820 => "0000000000000000", 18821 => "0000000000000000", 18822 => "0000000000000000", 18823 => "0000000000000000", 18824 => "0000000000000000", 18825 => "0000000000000000", 18826 => "0000000000000000", 18827 => "0000000000000000", 18828 => "0000000000000000", 18829 => "0000000000000000", 18830 => "0000000000000000", 18831 => "0000000000000000", 18832 => "0000000000000000", 18833 => "0000000000000000", 18834 => "0000000000000000", 18835 => "0000000000000000", 18836 => "0000000000000000", 18837 => "0000000000000000", 18838 => "0000000000000000", 18839 => "0000000000000000", 18840 => "0000000000000000", 18841 => "0000000000000000", 18842 => "0000000000000000", 18843 => "0000000000000000", 18844 => "0000000000000000", 18845 => "0000000000000000", 18846 => "0000000000000000", 18847 => "0000000000000000", 18848 => "0000000000000000", 18849 => "0000000000000000", 18850 => "0000000000000000", 18851 => "0000000000000000", 18852 => "0000000000000000", 18853 => "0000000000000000", 18854 => "0000000000000000", 18855 => "0000000000000000", 18856 => "0000000000000000", 18857 => "0000000000000000", 18858 => "0000000000000000", 18859 => "0000000000000000", 18860 => "0000000000000000", 18861 => "0000000000000000", 18862 => "0000000000000000", 18863 => "0000000000000000", 18864 => "0000000000000000", 18865 => "0000000000000000", 18866 => "0000000000000000", 18867 => "0000000000000000", 18868 => "0000000000000000", 18869 => "0000000000000000", 18870 => "0000000000000000", 18871 => "0000000000000000", 18872 => "0000000000000000", 18873 => "0000000000000000", 18874 => "0000000000000000", 18875 => "0000000000000000", 18876 => "0000000000000000", 18877 => "0000000000000000", 18878 => "0000000000000000", 18879 => "0000000000000000", 18880 => "0000000000000000", 18881 => "0000000000000000", 18882 => "0000000000000000", 18883 => "0000000000000000", 18884 => "0000000000000000", 18885 => "0000000000000000", 18886 => "0000000000000000", 18887 => "0000000000000000", 18888 => "0000000000000000", 18889 => "0000000000000000", 18890 => "0000000000000000", 18891 => "0000000000000000", 18892 => "0000000000000000", 18893 => "0000000000000000", 18894 => "0000000000000000", 18895 => "0000000000000000", 18896 => "0000000000000000", 18897 => "0000000000000000", 18898 => "0000000000000000", 18899 => "0000000000000000", 18900 => "0000000000000000", 18901 => "0000000000000000", 18902 => "0000000000000000", 18903 => "0000000000000000", 18904 => "0000000000000000", 18905 => "0000000000000000", 18906 => "0000000000000000", 18907 => "0000000000000000", 18908 => "0000000000000000", 18909 => "0000000000000000", 18910 => "0000000000000000", 18911 => "0000000000000000", 18912 => "0000000000000000", 18913 => "0000000000000000", 18914 => "0000000000000000", 18915 => "0000000000000000", 18916 => "0000000000000000", 18917 => "0000000000000000", 18918 => "0000000000000000", 18919 => "0000000000000000", 18920 => "0000000000000000", 18921 => "0000000000000000", 18922 => "0000000000000000", 18923 => "0000000000000000", 18924 => "0000000000000000", 18925 => "0000000000000000", 18926 => "0000000000000000", 18927 => "0000000000000000", 18928 => "0000000000000000", 18929 => "0000000000000000", 18930 => "0000000000000000", 18931 => "0000000000000000", 18932 => "0000000000000000", 18933 => "0000000000000000", 18934 => "0000000000000000", 18935 => "0000000000000000", 18936 => "0000000000000000", 18937 => "0000000000000000", 18938 => "0000000000000000", 18939 => "0000000000000000", 18940 => "0000000000000000", 18941 => "0000000000000000", 18942 => "0000000000000000", 18943 => "0000000000000000", 18944 => "0000000000000000", 18945 => "0000000000000000", 18946 => "0000000000000000", 18947 => "0000000000000000", 18948 => "0000000000000000", 18949 => "0000000000000000", 18950 => "0000000000000000", 18951 => "0000000000000000", 18952 => "0000000000000000", 18953 => "0000000000000000", 18954 => "0000000000000000", 18955 => "0000000000000000", 18956 => "0000000000000000", 18957 => "0000000000000000", 18958 => "0000000000000000", 18959 => "0000000000000000", 18960 => "0000000000000000", 18961 => "0000000000000000", 18962 => "0000000000000000", 18963 => "0000000000000000", 18964 => "0000000000000000", 18965 => "0000000000000000", 18966 => "0000000000000000", 18967 => "0000000000000000", 18968 => "0000000000000000", 18969 => "0000000000000000", 18970 => "0000000000000000", 18971 => "0000000000000000", 18972 => "0000000000000000", 18973 => "0000000000000000", 18974 => "0000000000000000", 18975 => "0000000000000000", 18976 => "0000000000000000", 18977 => "0000000000000000", 18978 => "0000000000000000", 18979 => "0000000000000000", 18980 => "0000000000000000", 18981 => "0000000000000000", 18982 => "0000000000000000", 18983 => "0000000000000000", 18984 => "0000000000000000", 18985 => "0000000000000000", 18986 => "0000000000000000", 18987 => "0000000000000000", 18988 => "0000000000000000", 18989 => "0000000000000000", 18990 => "0000000000000000", 18991 => "0000000000000000", 18992 => "0000000000000000", 18993 => "0000000000000000", 18994 => "0000000000000000", 18995 => "0000000000000000", 18996 => "0000000000000000", 18997 => "0000000000000000", 18998 => "0000000000000000", 18999 => "0000000000000000", 19000 => "0000000000000000", 19001 => "0000000000000000", 19002 => "0000000000000000", 19003 => "0000000000000000", 19004 => "0000000000000000", 19005 => "0000000000000000", 19006 => "0000000000000000", 19007 => "0000000000000000", 19008 => "0000000000000000", 19009 => "0000000000000000", 19010 => "0000000000000000", 19011 => "0000000000000000", 19012 => "0000000000000000", 19013 => "0000000000000000", 19014 => "0000000000000000", 19015 => "0000000000000000", 19016 => "0000000000000000", 19017 => "0000000000000000", 19018 => "0000000000000000", 19019 => "0000000000000000", 19020 => "0000000000000000", 19021 => "0000000000000000", 19022 => "0000000000000000", 19023 => "0000000000000000", 19024 => "0000000000000000", 19025 => "0000000000000000", 19026 => "0000000000000000", 19027 => "0000000000000000", 19028 => "0000000000000000", 19029 => "0000000000000000", 19030 => "0000000000000000", 19031 => "0000000000000000", 19032 => "0000000000000000", 19033 => "0000000000000000", 19034 => "0000000000000000", 19035 => "0000000000000000", 19036 => "0000000000000000", 19037 => "0000000000000000", 19038 => "0000000000000000", 19039 => "0000000000000000", 19040 => "0000000000000000", 19041 => "0000000000000000", 19042 => "0000000000000000", 19043 => "0000000000000000", 19044 => "0000000000000000", 19045 => "0000000000000000", 19046 => "0000000000000000", 19047 => "0000000000000000", 19048 => "0000000000000000", 19049 => "0000000000000000", 19050 => "0000000000000000", 19051 => "0000000000000000", 19052 => "0000000000000000", 19053 => "0000000000000000", 19054 => "0000000000000000", 19055 => "0000000000000000", 19056 => "0000000000000000", 19057 => "0000000000000000", 19058 => "0000000000000000", 19059 => "0000000000000000", 19060 => "0000000000000000", 19061 => "0000000000000000", 19062 => "0000000000000000", 19063 => "0000000000000000", 19064 => "0000000000000000", 19065 => "0000000000000000", 19066 => "0000000000000000", 19067 => "0000000000000000", 19068 => "0000000000000000", 19069 => "0000000000000000", 19070 => "0000000000000000", 19071 => "0000000000000000", 19072 => "0000000000000000", 19073 => "0000000000000000", 19074 => "0000000000000000", 19075 => "0000000000000000", 19076 => "0000000000000000", 19077 => "0000000000000000", 19078 => "0000000000000000", 19079 => "0000000000000000", 19080 => "0000000000000000", 19081 => "0000000000000000", 19082 => "0000000000000000", 19083 => "0000000000000000", 19084 => "0000000000000000", 19085 => "0000000000000000", 19086 => "0000000000000000", 19087 => "0000000000000000", 19088 => "0000000000000000", 19089 => "0000000000000000", 19090 => "0000000000000000", 19091 => "0000000000000000", 19092 => "0000000000000000", 19093 => "0000000000000000", 19094 => "0000000000000000", 19095 => "0000000000000000", 19096 => "0000000000000000", 19097 => "0000000000000000", 19098 => "0000000000000000", 19099 => "0000000000000000", 19100 => "0000000000000000", 19101 => "0000000000000000", 19102 => "0000000000000000", 19103 => "0000000000000000", 19104 => "0000000000000000", 19105 => "0000000000000000", 19106 => "0000000000000000", 19107 => "0000000000000000", 19108 => "0000000000000000", 19109 => "0000000000000000", 19110 => "0000000000000000", 19111 => "0000000000000000", 19112 => "0000000000000000", 19113 => "0000000000000000", 19114 => "0000000000000000", 19115 => "0000000000000000", 19116 => "0000000000000000", 19117 => "0000000000000000", 19118 => "0000000000000000", 19119 => "0000000000000000", 19120 => "0000000000000000", 19121 => "0000000000000000", 19122 => "0000000000000000", 19123 => "0000000000000000", 19124 => "0000000000000000", 19125 => "0000000000000000", 19126 => "0000000000000000", 19127 => "0000000000000000", 19128 => "0000000000000000", 19129 => "0000000000000000", 19130 => "0000000000000000", 19131 => "0000000000000000", 19132 => "0000000000000000", 19133 => "0000000000000000", 19134 => "0000000000000000", 19135 => "0000000000000000", 19136 => "0000000000000000", 19137 => "0000000000000000", 19138 => "0000000000000000", 19139 => "0000000000000000", 19140 => "0000000000000000", 19141 => "0000000000000000", 19142 => "0000000000000000", 19143 => "0000000000000000", 19144 => "0000000000000000", 19145 => "0000000000000000", 19146 => "0000000000000000", 19147 => "0000000000000000", 19148 => "0000000000000000", 19149 => "0000000000000000", 19150 => "0000000000000000", 19151 => "0000000000000000", 19152 => "0000000000000000", 19153 => "0000000000000000", 19154 => "0000000000000000", 19155 => "0000000000000000", 19156 => "0000000000000000", 19157 => "0000000000000000", 19158 => "0000000000000000", 19159 => "0000000000000000", 19160 => "0000000000000000", 19161 => "0000000000000000", 19162 => "0000000000000000", 19163 => "0000000000000000", 19164 => "0000000000000000", 19165 => "0000000000000000", 19166 => "0000000000000000", 19167 => "0000000000000000", 19168 => "0000000000000000", 19169 => "0000000000000000", 19170 => "0000000000000000", 19171 => "0000000000000000", 19172 => "0000000000000000", 19173 => "0000000000000000", 19174 => "0000000000000000", 19175 => "0000000000000000", 19176 => "0000000000000000", 19177 => "0000000000000000", 19178 => "0000000000000000", 19179 => "0000000000000000", 19180 => "0000000000000000", 19181 => "0000000000000000", 19182 => "0000000000000000", 19183 => "0000000000000000", 19184 => "0000000000000000", 19185 => "0000000000000000", 19186 => "0000000000000000", 19187 => "0000000000000000", 19188 => "0000000000000000", 19189 => "0000000000000000", 19190 => "0000000000000000", 19191 => "0000000000000000", 19192 => "0000000000000000", 19193 => "0000000000000000", 19194 => "0000000000000000", 19195 => "0000000000000000", 19196 => "0000000000000000", 19197 => "0000000000000000", 19198 => "0000000000000000", 19199 => "0000000000000000", 19200 => "0000000000000000", 19201 => "0000000000000000", 19202 => "0000000000000000", 19203 => "0000000000000000", 19204 => "0000000000000000", 19205 => "0000000000000000", 19206 => "0000000000000000", 19207 => "0000000000000000", 19208 => "0000000000000000", 19209 => "0000000000000000", 19210 => "0000000000000000", 19211 => "0000000000000000", 19212 => "0000000000000000", 19213 => "0000000000000000", 19214 => "0000000000000000", 19215 => "0000000000000000", 19216 => "0000000000000000", 19217 => "0000000000000000", 19218 => "0000000000000000", 19219 => "0000000000000000", 19220 => "0000000000000000", 19221 => "0000000000000000", 19222 => "0000000000000000", 19223 => "0000000000000000", 19224 => "0000000000000000", 19225 => "0000000000000000", 19226 => "0000000000000000", 19227 => "0000000000000000", 19228 => "0000000000000000", 19229 => "0000000000000000", 19230 => "0000000000000000", 19231 => "0000000000000000", 19232 => "0000000000000000", 19233 => "0000000000000000", 19234 => "0000000000000000", 19235 => "0000000000000000", 19236 => "0000000000000000", 19237 => "0000000000000000", 19238 => "0000000000000000", 19239 => "0000000000000000", 19240 => "0000000000000000", 19241 => "0000000000000000", 19242 => "0000000000000000", 19243 => "0000000000000000", 19244 => "0000000000000000", 19245 => "0000000000000000", 19246 => "0000000000000000", 19247 => "0000000000000000", 19248 => "0000000000000000", 19249 => "0000000000000000", 19250 => "0000000000000000", 19251 => "0000000000000000", 19252 => "0000000000000000", 19253 => "0000000000000000", 19254 => "0000000000000000", 19255 => "0000000000000000", 19256 => "0000000000000000", 19257 => "0000000000000000", 19258 => "0000000000000000", 19259 => "0000000000000000", 19260 => "0000000000000000", 19261 => "0000000000000000", 19262 => "0000000000000000", 19263 => "0000000000000000", 19264 => "0000000000000000", 19265 => "0000000000000000", 19266 => "0000000000000000", 19267 => "0000000000000000", 19268 => "0000000000000000", 19269 => "0000000000000000", 19270 => "0000000000000000", 19271 => "0000000000000000", 19272 => "0000000000000000", 19273 => "0000000000000000", 19274 => "0000000000000000", 19275 => "0000000000000000", 19276 => "0000000000000000", 19277 => "0000000000000000", 19278 => "0000000000000000", 19279 => "0000000000000000", 19280 => "0000000000000000", 19281 => "0000000000000000", 19282 => "0000000000000000", 19283 => "0000000000000000", 19284 => "0000000000000000", 19285 => "0000000000000000", 19286 => "0000000000000000", 19287 => "0000000000000000", 19288 => "0000000000000000", 19289 => "0000000000000000", 19290 => "0000000000000000", 19291 => "0000000000000000", 19292 => "0000000000000000", 19293 => "0000000000000000", 19294 => "0000000000000000", 19295 => "0000000000000000", 19296 => "0000000000000000", 19297 => "0000000000000000", 19298 => "0000000000000000", 19299 => "0000000000000000", 19300 => "0000000000000000", 19301 => "0000000000000000", 19302 => "0000000000000000", 19303 => "0000000000000000", 19304 => "0000000000000000", 19305 => "0000000000000000", 19306 => "0000000000000000", 19307 => "0000000000000000", 19308 => "0000000000000000", 19309 => "0000000000000000", 19310 => "0000000000000000", 19311 => "0000000000000000", 19312 => "0000000000000000", 19313 => "0000000000000000", 19314 => "0000000000000000", 19315 => "0000000000000000", 19316 => "0000000000000000", 19317 => "0000000000000000", 19318 => "0000000000000000", 19319 => "0000000000000000", 19320 => "0000000000000000", 19321 => "0000000000000000", 19322 => "0000000000000000", 19323 => "0000000000000000", 19324 => "0000000000000000", 19325 => "0000000000000000", 19326 => "0000000000000000", 19327 => "0000000000000000", 19328 => "0000000000000000", 19329 => "0000000000000000", 19330 => "0000000000000000", 19331 => "0000000000000000", 19332 => "0000000000000000", 19333 => "0000000000000000", 19334 => "0000000000000000", 19335 => "0000000000000000", 19336 => "0000000000000000", 19337 => "0000000000000000", 19338 => "0000000000000000", 19339 => "0000000000000000", 19340 => "0000000000000000", 19341 => "0000000000000000", 19342 => "0000000000000000", 19343 => "0000000000000000", 19344 => "0000000000000000", 19345 => "0000000000000000", 19346 => "0000000000000000", 19347 => "0000000000000000", 19348 => "0000000000000000", 19349 => "0000000000000000", 19350 => "0000000000000000", 19351 => "0000000000000000", 19352 => "0000000000000000", 19353 => "0000000000000000", 19354 => "0000000000000000", 19355 => "0000000000000000", 19356 => "0000000000000000", 19357 => "0000000000000000", 19358 => "0000000000000000", 19359 => "0000000000000000", 19360 => "0000000000000000", 19361 => "0000000000000000", 19362 => "0000000000000000", 19363 => "0000000000000000", 19364 => "0000000000000000", 19365 => "0000000000000000", 19366 => "0000000000000000", 19367 => "0000000000000000", 19368 => "0000000000000000", 19369 => "0000000000000000", 19370 => "0000000000000000", 19371 => "0000000000000000", 19372 => "0000000000000000", 19373 => "0000000000000000", 19374 => "0000000000000000", 19375 => "0000000000000000", 19376 => "0000000000000000", 19377 => "0000000000000000", 19378 => "0000000000000000", 19379 => "0000000000000000", 19380 => "0000000000000000", 19381 => "0000000000000000", 19382 => "0000000000000000", 19383 => "0000000000000000", 19384 => "0000000000000000", 19385 => "0000000000000000", 19386 => "0000000000000000", 19387 => "0000000000000000", 19388 => "0000000000000000", 19389 => "0000000000000000", 19390 => "0000000000000000", 19391 => "0000000000000000", 19392 => "0000000000000000", 19393 => "0000000000000000", 19394 => "0000000000000000", 19395 => "0000000000000000", 19396 => "0000000000000000", 19397 => "0000000000000000", 19398 => "0000000000000000", 19399 => "0000000000000000", 19400 => "0000000000000000", 19401 => "0000000000000000", 19402 => "0000000000000000", 19403 => "0000000000000000", 19404 => "0000000000000000", 19405 => "0000000000000000", 19406 => "0000000000000000", 19407 => "0000000000000000", 19408 => "0000000000000000", 19409 => "0000000000000000", 19410 => "0000000000000000", 19411 => "0000000000000000", 19412 => "0000000000000000", 19413 => "0000000000000000", 19414 => "0000000000000000", 19415 => "0000000000000000", 19416 => "0000000000000000", 19417 => "0000000000000000", 19418 => "0000000000000000", 19419 => "0000000000000000", 19420 => "0000000000000000", 19421 => "0000000000000000", 19422 => "0000000000000000", 19423 => "0000000000000000", 19424 => "0000000000000000", 19425 => "0000000000000000", 19426 => "0000000000000000", 19427 => "0000000000000000", 19428 => "0000000000000000", 19429 => "0000000000000000", 19430 => "0000000000000000", 19431 => "0000000000000000", 19432 => "0000000000000000", 19433 => "0000000000000000", 19434 => "0000000000000000", 19435 => "0000000000000000", 19436 => "0000000000000000", 19437 => "0000000000000000", 19438 => "0000000000000000", 19439 => "0000000000000000", 19440 => "0000000000000000", 19441 => "0000000000000000", 19442 => "0000000000000000", 19443 => "0000000000000000", 19444 => "0000000000000000", 19445 => "0000000000000000", 19446 => "0000000000000000", 19447 => "0000000000000000", 19448 => "0000000000000000", 19449 => "0000000000000000", 19450 => "0000000000000000", 19451 => "0000000000000000", 19452 => "0000000000000000", 19453 => "0000000000000000", 19454 => "0000000000000000", 19455 => "0000000000000000", 19456 => "0000000000000000", 19457 => "0000000000000000", 19458 => "0000000000000000", 19459 => "0000000000000000", 19460 => "0000000000000000", 19461 => "0000000000000000", 19462 => "0000000000000000", 19463 => "0000000000000000", 19464 => "0000000000000000", 19465 => "0000000000000000", 19466 => "0000000000000000", 19467 => "0000000000000000", 19468 => "0000000000000000", 19469 => "0000000000000000", 19470 => "0000000000000000", 19471 => "0000000000000000", 19472 => "0000000000000000", 19473 => "0000000000000000", 19474 => "0000000000000000", 19475 => "0000000000000000", 19476 => "0000000000000000", 19477 => "0000000000000000", 19478 => "0000000000000000", 19479 => "0000000000000000", 19480 => "0000000000000000", 19481 => "0000000000000000", 19482 => "0000000000000000", 19483 => "0000000000000000", 19484 => "0000000000000000", 19485 => "0000000000000000", 19486 => "0000000000000000", 19487 => "0000000000000000", 19488 => "0000000000000000", 19489 => "0000000000000000", 19490 => "0000000000000000", 19491 => "0000000000000000", 19492 => "0000000000000000", 19493 => "0000000000000000", 19494 => "0000000000000000", 19495 => "0000000000000000", 19496 => "0000000000000000", 19497 => "0000000000000000", 19498 => "0000000000000000", 19499 => "0000000000000000", 19500 => "0000000000000000", 19501 => "0000000000000000", 19502 => "0000000000000000", 19503 => "0000000000000000", 19504 => "0000000000000000", 19505 => "0000000000000000", 19506 => "0000000000000000", 19507 => "0000000000000000", 19508 => "0000000000000000", 19509 => "0000000000000000", 19510 => "0000000000000000", 19511 => "0000000000000000", 19512 => "0000000000000000", 19513 => "0000000000000000", 19514 => "0000000000000000", 19515 => "0000000000000000", 19516 => "0000000000000000", 19517 => "0000000000000000", 19518 => "0000000000000000", 19519 => "0000000000000000", 19520 => "0000000000000000", 19521 => "0000000000000000", 19522 => "0000000000000000", 19523 => "0000000000000000", 19524 => "0000000000000000", 19525 => "0000000000000000", 19526 => "0000000000000000", 19527 => "0000000000000000", 19528 => "0000000000000000", 19529 => "0000000000000000", 19530 => "0000000000000000", 19531 => "0000000000000000", 19532 => "0000000000000000", 19533 => "0000000000000000", 19534 => "0000000000000000", 19535 => "0000000000000000", 19536 => "0000000000000000", 19537 => "0000000000000000", 19538 => "0000000000000000", 19539 => "0000000000000000", 19540 => "0000000000000000", 19541 => "0000000000000000", 19542 => "0000000000000000", 19543 => "0000000000000000", 19544 => "0000000000000000", 19545 => "0000000000000000", 19546 => "0000000000000000", 19547 => "0000000000000000", 19548 => "0000000000000000", 19549 => "0000000000000000", 19550 => "0000000000000000", 19551 => "0000000000000000", 19552 => "0000000000000000", 19553 => "0000000000000000", 19554 => "0000000000000000", 19555 => "0000000000000000", 19556 => "0000000000000000", 19557 => "0000000000000000", 19558 => "0000000000000000", 19559 => "0000000000000000", 19560 => "0000000000000000", 19561 => "0000000000000000", 19562 => "0000000000000000", 19563 => "0000000000000000", 19564 => "0000000000000000", 19565 => "0000000000000000", 19566 => "0000000000000000", 19567 => "0000000000000000", 19568 => "0000000000000000", 19569 => "0000000000000000", 19570 => "0000000000000000", 19571 => "0000000000000000", 19572 => "0000000000000000", 19573 => "0000000000000000", 19574 => "0000000000000000", 19575 => "0000000000000000", 19576 => "0000000000000000", 19577 => "0000000000000000", 19578 => "0000000000000000", 19579 => "0000000000000000", 19580 => "0000000000000000", 19581 => "0000000000000000", 19582 => "0000000000000000", 19583 => "0000000000000000", 19584 => "0000000000000000", 19585 => "0000000000000000", 19586 => "0000000000000000", 19587 => "0000000000000000", 19588 => "0000000000000000", 19589 => "0000000000000000", 19590 => "0000000000000000", 19591 => "0000000000000000", 19592 => "0000000000000000", 19593 => "0000000000000000", 19594 => "0000000000000000", 19595 => "0000000000000000", 19596 => "0000000000000000", 19597 => "0000000000000000", 19598 => "0000000000000000", 19599 => "0000000000000000", 19600 => "0000000000000000", 19601 => "0000000000000000", 19602 => "0000000000000000", 19603 => "0000000000000000", 19604 => "0000000000000000", 19605 => "0000000000000000", 19606 => "0000000000000000", 19607 => "0000000000000000", 19608 => "0000000000000000", 19609 => "0000000000000000", 19610 => "0000000000000000", 19611 => "0000000000000000", 19612 => "0000000000000000", 19613 => "0000000000000000", 19614 => "0000000000000000", 19615 => "0000000000000000", 19616 => "0000000000000000", 19617 => "0000000000000000", 19618 => "0000000000000000", 19619 => "0000000000000000", 19620 => "0000000000000000", 19621 => "0000000000000000", 19622 => "0000000000000000", 19623 => "0000000000000000", 19624 => "0000000000000000", 19625 => "0000000000000000", 19626 => "0000000000000000", 19627 => "0000000000000000", 19628 => "0000000000000000", 19629 => "0000000000000000", 19630 => "0000000000000000", 19631 => "0000000000000000", 19632 => "0000000000000000", 19633 => "0000000000000000", 19634 => "0000000000000000", 19635 => "0000000000000000", 19636 => "0000000000000000", 19637 => "0000000000000000", 19638 => "0000000000000000", 19639 => "0000000000000000", 19640 => "0000000000000000", 19641 => "0000000000000000", 19642 => "0000000000000000", 19643 => "0000000000000000", 19644 => "0000000000000000", 19645 => "0000000000000000", 19646 => "0000000000000000", 19647 => "0000000000000000", 19648 => "0000000000000000", 19649 => "0000000000000000", 19650 => "0000000000000000", 19651 => "0000000000000000", 19652 => "0000000000000000", 19653 => "0000000000000000", 19654 => "0000000000000000", 19655 => "0000000000000000", 19656 => "0000000000000000", 19657 => "0000000000000000", 19658 => "0000000000000000", 19659 => "0000000000000000", 19660 => "0000000000000000", 19661 => "0000000000000000", 19662 => "0000000000000000", 19663 => "0000000000000000", 19664 => "0000000000000000", 19665 => "0000000000000000", 19666 => "0000000000000000", 19667 => "0000000000000000", 19668 => "0000000000000000", 19669 => "0000000000000000", 19670 => "0000000000000000", 19671 => "0000000000000000", 19672 => "0000000000000000", 19673 => "0000000000000000", 19674 => "0000000000000000", 19675 => "0000000000000000", 19676 => "0000000000000000", 19677 => "0000000000000000", 19678 => "0000000000000000", 19679 => "0000000000000000", 19680 => "0000000000000000", 19681 => "0000000000000000", 19682 => "0000000000000000", 19683 => "0000000000000000", 19684 => "0000000000000000", 19685 => "0000000000000000", 19686 => "0000000000000000", 19687 => "0000000000000000", 19688 => "0000000000000000", 19689 => "0000000000000000", 19690 => "0000000000000000", 19691 => "0000000000000000", 19692 => "0000000000000000", 19693 => "0000000000000000", 19694 => "0000000000000000", 19695 => "0000000000000000", 19696 => "0000000000000000", 19697 => "0000000000000000", 19698 => "0000000000000000", 19699 => "0000000000000000", 19700 => "0000000000000000", 19701 => "0000000000000000", 19702 => "0000000000000000", 19703 => "0000000000000000", 19704 => "0000000000000000", 19705 => "0000000000000000", 19706 => "0000000000000000", 19707 => "0000000000000000", 19708 => "0000000000000000", 19709 => "0000000000000000", 19710 => "0000000000000000", 19711 => "0000000000000000", 19712 => "0000000000000000", 19713 => "0000000000000000", 19714 => "0000000000000000", 19715 => "0000000000000000", 19716 => "0000000000000000", 19717 => "0000000000000000", 19718 => "0000000000000000", 19719 => "0000000000000000", 19720 => "0000000000000000", 19721 => "0000000000000000", 19722 => "0000000000000000", 19723 => "0000000000000000", 19724 => "0000000000000000", 19725 => "0000000000000000", 19726 => "0000000000000000", 19727 => "0000000000000000", 19728 => "0000000000000000", 19729 => "0000000000000000", 19730 => "0000000000000000", 19731 => "0000000000000000", 19732 => "0000000000000000", 19733 => "0000000000000000", 19734 => "0000000000000000", 19735 => "0000000000000000", 19736 => "0000000000000000", 19737 => "0000000000000000", 19738 => "0000000000000000", 19739 => "0000000000000000", 19740 => "0000000000000000", 19741 => "0000000000000000", 19742 => "0000000000000000", 19743 => "0000000000000000", 19744 => "0000000000000000", 19745 => "0000000000000000", 19746 => "0000000000000000", 19747 => "0000000000000000", 19748 => "0000000000000000", 19749 => "0000000000000000", 19750 => "0000000000000000", 19751 => "0000000000000000", 19752 => "0000000000000000", 19753 => "0000000000000000", 19754 => "0000000000000000", 19755 => "0000000000000000", 19756 => "0000000000000000", 19757 => "0000000000000000", 19758 => "0000000000000000", 19759 => "0000000000000000", 19760 => "0000000000000000", 19761 => "0000000000000000", 19762 => "0000000000000000", 19763 => "0000000000000000", 19764 => "0000000000000000", 19765 => "0000000000000000", 19766 => "0000000000000000", 19767 => "0000000000000000", 19768 => "0000000000000000", 19769 => "0000000000000000", 19770 => "0000000000000000", 19771 => "0000000000000000", 19772 => "0000000000000000", 19773 => "0000000000000000", 19774 => "0000000000000000", 19775 => "0000000000000000", 19776 => "0000000000000000", 19777 => "0000000000000000", 19778 => "0000000000000000", 19779 => "0000000000000000", 19780 => "0000000000000000", 19781 => "0000000000000000", 19782 => "0000000000000000", 19783 => "0000000000000000", 19784 => "0000000000000000", 19785 => "0000000000000000", 19786 => "0000000000000000", 19787 => "0000000000000000", 19788 => "0000000000000000", 19789 => "0000000000000000", 19790 => "0000000000000000", 19791 => "0000000000000000", 19792 => "0000000000000000", 19793 => "0000000000000000", 19794 => "0000000000000000", 19795 => "0000000000000000", 19796 => "0000000000000000", 19797 => "0000000000000000", 19798 => "0000000000000000", 19799 => "0000000000000000", 19800 => "0000000000000000", 19801 => "0000000000000000", 19802 => "0000000000000000", 19803 => "0000000000000000", 19804 => "0000000000000000", 19805 => "0000000000000000", 19806 => "0000000000000000", 19807 => "0000000000000000", 19808 => "0000000000000000", 19809 => "0000000000000000", 19810 => "0000000000000000", 19811 => "0000000000000000", 19812 => "0000000000000000", 19813 => "0000000000000000", 19814 => "0000000000000000", 19815 => "0000000000000000", 19816 => "0000000000000000", 19817 => "0000000000000000", 19818 => "0000000000000000", 19819 => "0000000000000000", 19820 => "0000000000000000", 19821 => "0000000000000000", 19822 => "0000000000000000", 19823 => "0000000000000000", 19824 => "0000000000000000", 19825 => "0000000000000000", 19826 => "0000000000000000", 19827 => "0000000000000000", 19828 => "0000000000000000", 19829 => "0000000000000000", 19830 => "0000000000000000", 19831 => "0000000000000000", 19832 => "0000000000000000", 19833 => "0000000000000000", 19834 => "0000000000000000", 19835 => "0000000000000000", 19836 => "0000000000000000", 19837 => "0000000000000000", 19838 => "0000000000000000", 19839 => "0000000000000000", 19840 => "0000000000000000", 19841 => "0000000000000000", 19842 => "0000000000000000", 19843 => "0000000000000000", 19844 => "0000000000000000", 19845 => "0000000000000000", 19846 => "0000000000000000", 19847 => "0000000000000000", 19848 => "0000000000000000", 19849 => "0000000000000000", 19850 => "0000000000000000", 19851 => "0000000000000000", 19852 => "0000000000000000", 19853 => "0000000000000000", 19854 => "0000000000000000", 19855 => "0000000000000000", 19856 => "0000000000000000", 19857 => "0000000000000000", 19858 => "0000000000000000", 19859 => "0000000000000000", 19860 => "0000000000000000", 19861 => "0000000000000000", 19862 => "0000000000000000", 19863 => "0000000000000000", 19864 => "0000000000000000", 19865 => "0000000000000000", 19866 => "0000000000000000", 19867 => "0000000000000000", 19868 => "0000000000000000", 19869 => "0000000000000000", 19870 => "0000000000000000", 19871 => "0000000000000000", 19872 => "0000000000000000", 19873 => "0000000000000000", 19874 => "0000000000000000", 19875 => "0000000000000000", 19876 => "0000000000000000", 19877 => "0000000000000000", 19878 => "0000000000000000", 19879 => "0000000000000000", 19880 => "0000000000000000", 19881 => "0000000000000000", 19882 => "0000000000000000", 19883 => "0000000000000000", 19884 => "0000000000000000", 19885 => "0000000000000000", 19886 => "0000000000000000", 19887 => "0000000000000000", 19888 => "0000000000000000", 19889 => "0000000000000000", 19890 => "0000000000000000", 19891 => "0000000000000000", 19892 => "0000000000000000", 19893 => "0000000000000000", 19894 => "0000000000000000", 19895 => "0000000000000000", 19896 => "0000000000000000", 19897 => "0000000000000000", 19898 => "0000000000000000", 19899 => "0000000000000000", 19900 => "0000000000000000", 19901 => "0000000000000000", 19902 => "0000000000000000", 19903 => "0000000000000000", 19904 => "0000000000000000", 19905 => "0000000000000000", 19906 => "0000000000000000", 19907 => "0000000000000000", 19908 => "0000000000000000", 19909 => "0000000000000000", 19910 => "0000000000000000", 19911 => "0000000000000000", 19912 => "0000000000000000", 19913 => "0000000000000000", 19914 => "0000000000000000", 19915 => "0000000000000000", 19916 => "0000000000000000", 19917 => "0000000000000000", 19918 => "0000000000000000", 19919 => "0000000000000000", 19920 => "0000000000000000", 19921 => "0000000000000000", 19922 => "0000000000000000", 19923 => "0000000000000000", 19924 => "0000000000000000", 19925 => "0000000000000000", 19926 => "0000000000000000", 19927 => "0000000000000000", 19928 => "0000000000000000", 19929 => "0000000000000000", 19930 => "0000000000000000", 19931 => "0000000000000000", 19932 => "0000000000000000", 19933 => "0000000000000000", 19934 => "0000000000000000", 19935 => "0000000000000000", 19936 => "0000000000000000", 19937 => "0000000000000000", 19938 => "0000000000000000", 19939 => "0000000000000000", 19940 => "0000000000000000", 19941 => "0000000000000000", 19942 => "0000000000000000", 19943 => "0000000000000000", 19944 => "0000000000000000", 19945 => "0000000000000000", 19946 => "0000000000000000", 19947 => "0000000000000000", 19948 => "0000000000000000", 19949 => "0000000000000000", 19950 => "0000000000000000", 19951 => "0000000000000000", 19952 => "0000000000000000", 19953 => "0000000000000000", 19954 => "0000000000000000", 19955 => "0000000000000000", 19956 => "0000000000000000", 19957 => "0000000000000000", 19958 => "0000000000000000", 19959 => "0000000000000000", 19960 => "0000000000000000", 19961 => "0000000000000000", 19962 => "0000000000000000", 19963 => "0000000000000000", 19964 => "0000000000000000", 19965 => "0000000000000000", 19966 => "0000000000000000", 19967 => "0000000000000000", 19968 => "0000000000000000", 19969 => "0000000000000000", 19970 => "0000000000000000", 19971 => "0000000000000000", 19972 => "0000000000000000", 19973 => "0000000000000000", 19974 => "0000000000000000", 19975 => "0000000000000000", 19976 => "0000000000000000", 19977 => "0000000000000000", 19978 => "0000000000000000", 19979 => "0000000000000000", 19980 => "0000000000000000", 19981 => "0000000000000000", 19982 => "0000000000000000", 19983 => "0000000000000000", 19984 => "0000000000000000", 19985 => "0000000000000000", 19986 => "0000000000000000", 19987 => "0000000000000000", 19988 => "0000000000000000", 19989 => "0000000000000000", 19990 => "0000000000000000", 19991 => "0000000000000000", 19992 => "0000000000000000", 19993 => "0000000000000000", 19994 => "0000000000000000", 19995 => "0000000000000000", 19996 => "0000000000000000", 19997 => "0000000000000000", 19998 => "0000000000000000", 19999 => "0000000000000000", 20000 => "0000000000000000", 20001 => "0000000000000000", 20002 => "0000000000000000", 20003 => "0000000000000000", 20004 => "0000000000000000", 20005 => "0000000000000000", 20006 => "0000000000000000", 20007 => "0000000000000000", 20008 => "0000000000000000", 20009 => "0000000000000000", 20010 => "0000000000000000", 20011 => "0000000000000000", 20012 => "0000000000000000", 20013 => "0000000000000000", 20014 => "0000000000000000", 20015 => "0000000000000000", 20016 => "0000000000000000", 20017 => "0000000000000000", 20018 => "0000000000000000", 20019 => "0000000000000000", 20020 => "0000000000000000", 20021 => "0000000000000000", 20022 => "0000000000000000", 20023 => "0000000000000000", 20024 => "0000000000000000", 20025 => "0000000000000000", 20026 => "0000000000000000", 20027 => "0000000000000000", 20028 => "0000000000000000", 20029 => "0000000000000000", 20030 => "0000000000000000", 20031 => "0000000000000000", 20032 => "0000000000000000", 20033 => "0000000000000000", 20034 => "0000000000000000", 20035 => "0000000000000000", 20036 => "0000000000000000", 20037 => "0000000000000000", 20038 => "0000000000000000", 20039 => "0000000000000000", 20040 => "0000000000000000", 20041 => "0000000000000000", 20042 => "0000000000000000", 20043 => "0000000000000000", 20044 => "0000000000000000", 20045 => "0000000000000000", 20046 => "0000000000000000", 20047 => "0000000000000000", 20048 => "0000000000000000", 20049 => "0000000000000000", 20050 => "0000000000000000", 20051 => "0000000000000000", 20052 => "0000000000000000", 20053 => "0000000000000000", 20054 => "0000000000000000", 20055 => "0000000000000000", 20056 => "0000000000000000", 20057 => "0000000000000000", 20058 => "0000000000000000", 20059 => "0000000000000000", 20060 => "0000000000000000", 20061 => "0000000000000000", 20062 => "0000000000000000", 20063 => "0000000000000000", 20064 => "0000000000000000", 20065 => "0000000000000000", 20066 => "0000000000000000", 20067 => "0000000000000000", 20068 => "0000000000000000", 20069 => "0000000000000000", 20070 => "0000000000000000", 20071 => "0000000000000000", 20072 => "0000000000000000", 20073 => "0000000000000000", 20074 => "0000000000000000", 20075 => "0000000000000000", 20076 => "0000000000000000", 20077 => "0000000000000000", 20078 => "0000000000000000", 20079 => "0000000000000000", 20080 => "0000000000000000", 20081 => "0000000000000000", 20082 => "0000000000000000", 20083 => "0000000000000000", 20084 => "0000000000000000", 20085 => "0000000000000000", 20086 => "0000000000000000", 20087 => "0000000000000000", 20088 => "0000000000000000", 20089 => "0000000000000000", 20090 => "0000000000000000", 20091 => "0000000000000000", 20092 => "0000000000000000", 20093 => "0000000000000000", 20094 => "0000000000000000", 20095 => "0000000000000000", 20096 => "0000000000000000", 20097 => "0000000000000000", 20098 => "0000000000000000", 20099 => "0000000000000000", 20100 => "0000000000000000", 20101 => "0000000000000000", 20102 => "0000000000000000", 20103 => "0000000000000000", 20104 => "0000000000000000", 20105 => "0000000000000000", 20106 => "0000000000000000", 20107 => "0000000000000000", 20108 => "0000000000000000", 20109 => "0000000000000000", 20110 => "0000000000000000", 20111 => "0000000000000000", 20112 => "0000000000000000", 20113 => "0000000000000000", 20114 => "0000000000000000", 20115 => "0000000000000000", 20116 => "0000000000000000", 20117 => "0000000000000000", 20118 => "0000000000000000", 20119 => "0000000000000000", 20120 => "0000000000000000", 20121 => "0000000000000000", 20122 => "0000000000000000", 20123 => "0000000000000000", 20124 => "0000000000000000", 20125 => "0000000000000000", 20126 => "0000000000000000", 20127 => "0000000000000000", 20128 => "0000000000000000", 20129 => "0000000000000000", 20130 => "0000000000000000", 20131 => "0000000000000000", 20132 => "0000000000000000", 20133 => "0000000000000000", 20134 => "0000000000000000", 20135 => "0000000000000000", 20136 => "0000000000000000", 20137 => "0000000000000000", 20138 => "0000000000000000", 20139 => "0000000000000000", 20140 => "0000000000000000", 20141 => "0000000000000000", 20142 => "0000000000000000", 20143 => "0000000000000000", 20144 => "0000000000000000", 20145 => "0000000000000000", 20146 => "0000000000000000", 20147 => "0000000000000000", 20148 => "0000000000000000", 20149 => "0000000000000000", 20150 => "0000000000000000", 20151 => "0000000000000000", 20152 => "0000000000000000", 20153 => "0000000000000000", 20154 => "0000000000000000", 20155 => "0000000000000000", 20156 => "0000000000000000", 20157 => "0000000000000000", 20158 => "0000000000000000", 20159 => "0000000000000000", 20160 => "0000000000000000", 20161 => "0000000000000000", 20162 => "0000000000000000", 20163 => "0000000000000000", 20164 => "0000000000000000", 20165 => "0000000000000000", 20166 => "0000000000000000", 20167 => "0000000000000000", 20168 => "0000000000000000", 20169 => "0000000000000000", 20170 => "0000000000000000", 20171 => "0000000000000000", 20172 => "0000000000000000", 20173 => "0000000000000000", 20174 => "0000000000000000", 20175 => "0000000000000000", 20176 => "0000000000000000", 20177 => "0000000000000000", 20178 => "0000000000000000", 20179 => "0000000000000000", 20180 => "0000000000000000", 20181 => "0000000000000000", 20182 => "0000000000000000", 20183 => "0000000000000000", 20184 => "0000000000000000", 20185 => "0000000000000000", 20186 => "0000000000000000", 20187 => "0000000000000000", 20188 => "0000000000000000", 20189 => "0000000000000000", 20190 => "0000000000000000", 20191 => "0000000000000000", 20192 => "0000000000000000", 20193 => "0000000000000000", 20194 => "0000000000000000", 20195 => "0000000000000000", 20196 => "0000000000000000", 20197 => "0000000000000000", 20198 => "0000000000000000", 20199 => "0000000000000000", 20200 => "0000000000000000", 20201 => "0000000000000000", 20202 => "0000000000000000", 20203 => "0000000000000000", 20204 => "0000000000000000", 20205 => "0000000000000000", 20206 => "0000000000000000", 20207 => "0000000000000000", 20208 => "0000000000000000", 20209 => "0000000000000000", 20210 => "0000000000000000", 20211 => "0000000000000000", 20212 => "0000000000000000", 20213 => "0000000000000000", 20214 => "0000000000000000", 20215 => "0000000000000000", 20216 => "0000000000000000", 20217 => "0000000000000000", 20218 => "0000000000000000", 20219 => "0000000000000000", 20220 => "0000000000000000", 20221 => "0000000000000000", 20222 => "0000000000000000", 20223 => "0000000000000000", 20224 => "0000000000000000", 20225 => "0000000000000000", 20226 => "0000000000000000", 20227 => "0000000000000000", 20228 => "0000000000000000", 20229 => "0000000000000000", 20230 => "0000000000000000", 20231 => "0000000000000000", 20232 => "0000000000000000", 20233 => "0000000000000000", 20234 => "0000000000000000", 20235 => "0000000000000000", 20236 => "0000000000000000", 20237 => "0000000000000000", 20238 => "0000000000000000", 20239 => "0000000000000000", 20240 => "0000000000000000", 20241 => "0000000000000000", 20242 => "0000000000000000", 20243 => "0000000000000000", 20244 => "0000000000000000", 20245 => "0000000000000000", 20246 => "0000000000000000", 20247 => "0000000000000000", 20248 => "0000000000000000", 20249 => "0000000000000000", 20250 => "0000000000000000", 20251 => "0000000000000000", 20252 => "0000000000000000", 20253 => "0000000000000000", 20254 => "0000000000000000", 20255 => "0000000000000000", 20256 => "0000000000000000", 20257 => "0000000000000000", 20258 => "0000000000000000", 20259 => "0000000000000000", 20260 => "0000000000000000", 20261 => "0000000000000000", 20262 => "0000000000000000", 20263 => "0000000000000000", 20264 => "0000000000000000", 20265 => "0000000000000000", 20266 => "0000000000000000", 20267 => "0000000000000000", 20268 => "0000000000000000", 20269 => "0000000000000000", 20270 => "0000000000000000", 20271 => "0000000000000000", 20272 => "0000000000000000", 20273 => "0000000000000000", 20274 => "0000000000000000", 20275 => "0000000000000000", 20276 => "0000000000000000", 20277 => "0000000000000000", 20278 => "0000000000000000", 20279 => "0000000000000000", 20280 => "0000000000000000", 20281 => "0000000000000000", 20282 => "0000000000000000", 20283 => "0000000000000000", 20284 => "0000000000000000", 20285 => "0000000000000000", 20286 => "0000000000000000", 20287 => "0000000000000000", 20288 => "0000000000000000", 20289 => "0000000000000000", 20290 => "0000000000000000", 20291 => "0000000000000000", 20292 => "0000000000000000", 20293 => "0000000000000000", 20294 => "0000000000000000", 20295 => "0000000000000000", 20296 => "0000000000000000", 20297 => "0000000000000000", 20298 => "0000000000000000", 20299 => "0000000000000000", 20300 => "0000000000000000", 20301 => "0000000000000000", 20302 => "0000000000000000", 20303 => "0000000000000000", 20304 => "0000000000000000", 20305 => "0000000000000000", 20306 => "0000000000000000", 20307 => "0000000000000000", 20308 => "0000000000000000", 20309 => "0000000000000000", 20310 => "0000000000000000", 20311 => "0000000000000000", 20312 => "0000000000000000", 20313 => "0000000000000000", 20314 => "0000000000000000", 20315 => "0000000000000000", 20316 => "0000000000000000", 20317 => "0000000000000000", 20318 => "0000000000000000", 20319 => "0000000000000000", 20320 => "0000000000000000", 20321 => "0000000000000000", 20322 => "0000000000000000", 20323 => "0000000000000000", 20324 => "0000000000000000", 20325 => "0000000000000000", 20326 => "0000000000000000", 20327 => "0000000000000000", 20328 => "0000000000000000", 20329 => "0000000000000000", 20330 => "0000000000000000", 20331 => "0000000000000000", 20332 => "0000000000000000", 20333 => "0000000000000000", 20334 => "0000000000000000", 20335 => "0000000000000000", 20336 => "0000000000000000", 20337 => "0000000000000000", 20338 => "0000000000000000", 20339 => "0000000000000000", 20340 => "0000000000000000", 20341 => "0000000000000000", 20342 => "0000000000000000", 20343 => "0000000000000000", 20344 => "0000000000000000", 20345 => "0000000000000000", 20346 => "0000000000000000", 20347 => "0000000000000000", 20348 => "0000000000000000", 20349 => "0000000000000000", 20350 => "0000000000000000", 20351 => "0000000000000000", 20352 => "0000000000000000", 20353 => "0000000000000000", 20354 => "0000000000000000", 20355 => "0000000000000000", 20356 => "0000000000000000", 20357 => "0000000000000000", 20358 => "0000000000000000", 20359 => "0000000000000000", 20360 => "0000000000000000", 20361 => "0000000000000000", 20362 => "0000000000000000", 20363 => "0000000000000000", 20364 => "0000000000000000", 20365 => "0000000000000000", 20366 => "0000000000000000", 20367 => "0000000000000000", 20368 => "0000000000000000", 20369 => "0000000000000000", 20370 => "0000000000000000", 20371 => "0000000000000000", 20372 => "0000000000000000", 20373 => "0000000000000000", 20374 => "0000000000000000", 20375 => "0000000000000000", 20376 => "0000000000000000", 20377 => "0000000000000000", 20378 => "0000000000000000", 20379 => "0000000000000000", 20380 => "0000000000000000", 20381 => "0000000000000000", 20382 => "0000000000000000", 20383 => "0000000000000000", 20384 => "0000000000000000", 20385 => "0000000000000000", 20386 => "0000000000000000", 20387 => "0000000000000000", 20388 => "0000000000000000", 20389 => "0000000000000000", 20390 => "0000000000000000", 20391 => "0000000000000000", 20392 => "0000000000000000", 20393 => "0000000000000000", 20394 => "0000000000000000", 20395 => "0000000000000000", 20396 => "0000000000000000", 20397 => "0000000000000000", 20398 => "0000000000000000", 20399 => "0000000000000000", 20400 => "0000000000000000", 20401 => "0000000000000000", 20402 => "0000000000000000", 20403 => "0000000000000000", 20404 => "0000000000000000", 20405 => "0000000000000000", 20406 => "0000000000000000", 20407 => "0000000000000000", 20408 => "0000000000000000", 20409 => "0000000000000000", 20410 => "0000000000000000", 20411 => "0000000000000000", 20412 => "0000000000000000", 20413 => "0000000000000000", 20414 => "0000000000000000", 20415 => "0000000000000000", 20416 => "0000000000000000", 20417 => "0000000000000000", 20418 => "0000000000000000", 20419 => "0000000000000000", 20420 => "0000000000000000", 20421 => "0000000000000000", 20422 => "0000000000000000", 20423 => "0000000000000000", 20424 => "0000000000000000", 20425 => "0000000000000000", 20426 => "0000000000000000", 20427 => "0000000000000000", 20428 => "0000000000000000", 20429 => "0000000000000000", 20430 => "0000000000000000", 20431 => "0000000000000000", 20432 => "0000000000000000", 20433 => "0000000000000000", 20434 => "0000000000000000", 20435 => "0000000000000000", 20436 => "0000000000000000", 20437 => "0000000000000000", 20438 => "0000000000000000", 20439 => "0000000000000000", 20440 => "0000000000000000", 20441 => "0000000000000000", 20442 => "0000000000000000", 20443 => "0000000000000000", 20444 => "0000000000000000", 20445 => "0000000000000000", 20446 => "0000000000000000", 20447 => "0000000000000000", 20448 => "0000000000000000", 20449 => "0000000000000000", 20450 => "0000000000000000", 20451 => "0000000000000000", 20452 => "0000000000000000", 20453 => "0000000000000000", 20454 => "0000000000000000", 20455 => "0000000000000000", 20456 => "0000000000000000", 20457 => "0000000000000000", 20458 => "0000000000000000", 20459 => "0000000000000000", 20460 => "0000000000000000", 20461 => "0000000000000000", 20462 => "0000000000000000", 20463 => "0000000000000000", 20464 => "0000000000000000", 20465 => "0000000000000000", 20466 => "0000000000000000", 20467 => "0000000000000000", 20468 => "0000000000000000", 20469 => "0000000000000000", 20470 => "0000000000000000", 20471 => "0000000000000000", 20472 => "0000000000000000", 20473 => "0000000000000000", 20474 => "0000000000000000", 20475 => "0000000000000000", 20476 => "0000000000000000", 20477 => "0000000000000000", 20478 => "0000000000000000", 20479 => "0000000000000000", 20480 => "0000000000000000", 20481 => "0000000000000000", 20482 => "0000000000000000", 20483 => "0000000000000000", 20484 => "0000000000000000", 20485 => "0000000000000000", 20486 => "0000000000000000", 20487 => "0000000000000000", 20488 => "0000000000000000", 20489 => "0000000000000000", 20490 => "0000000000000000", 20491 => "0000000000000000", 20492 => "0000000000000000", 20493 => "0000000000000000", 20494 => "0000000000000000", 20495 => "0000000000000000", 20496 => "0000000000000000", 20497 => "0000000000000000", 20498 => "0000000000000000", 20499 => "0000000000000000", 20500 => "0000000000000000", 20501 => "0000000000000000", 20502 => "0000000000000000", 20503 => "0000000000000000", 20504 => "0000000000000000", 20505 => "0000000000000000", 20506 => "0000000000000000", 20507 => "0000000000000000", 20508 => "0000000000000000", 20509 => "0000000000000000", 20510 => "0000000000000000", 20511 => "0000000000000000", 20512 => "0000000000000000", 20513 => "0000000000000000", 20514 => "0000000000000000", 20515 => "0000000000000000", 20516 => "0000000000000000", 20517 => "0000000000000000", 20518 => "0000000000000000", 20519 => "0000000000000000", 20520 => "0000000000000000", 20521 => "0000000000000000", 20522 => "0000000000000000", 20523 => "0000000000000000", 20524 => "0000000000000000", 20525 => "0000000000000000", 20526 => "0000000000000000", 20527 => "0000000000000000", 20528 => "0000000000000000", 20529 => "0000000000000000", 20530 => "0000000000000000", 20531 => "0000000000000000", 20532 => "0000000000000000", 20533 => "0000000000000000", 20534 => "0000000000000000", 20535 => "0000000000000000", 20536 => "0000000000000000", 20537 => "0000000000000000", 20538 => "0000000000000000", 20539 => "0000000000000000", 20540 => "0000000000000000", 20541 => "0000000000000000", 20542 => "0000000000000000", 20543 => "0000000000000000", 20544 => "0000000000000000", 20545 => "0000000000000000", 20546 => "0000000000000000", 20547 => "0000000000000000", 20548 => "0000000000000000", 20549 => "0000000000000000", 20550 => "0000000000000000", 20551 => "0000000000000000", 20552 => "0000000000000000", 20553 => "0000000000000000", 20554 => "0000000000000000", 20555 => "0000000000000000", 20556 => "0000000000000000", 20557 => "0000000000000000", 20558 => "0000000000000000", 20559 => "0000000000000000", 20560 => "0000000000000000", 20561 => "0000000000000000", 20562 => "0000000000000000", 20563 => "0000000000000000", 20564 => "0000000000000000", 20565 => "0000000000000000", 20566 => "0000000000000000", 20567 => "0000000000000000", 20568 => "0000000000000000", 20569 => "0000000000000000", 20570 => "0000000000000000", 20571 => "0000000000000000", 20572 => "0000000000000000", 20573 => "0000000000000000", 20574 => "0000000000000000", 20575 => "0000000000000000", 20576 => "0000000000000000", 20577 => "0000000000000000", 20578 => "0000000000000000", 20579 => "0000000000000000", 20580 => "0000000000000000", 20581 => "0000000000000000", 20582 => "0000000000000000", 20583 => "0000000000000000", 20584 => "0000000000000000", 20585 => "0000000000000000", 20586 => "0000000000000000", 20587 => "0000000000000000", 20588 => "0000000000000000", 20589 => "0000000000000000", 20590 => "0000000000000000", 20591 => "0000000000000000", 20592 => "0000000000000000", 20593 => "0000000000000000", 20594 => "0000000000000000", 20595 => "0000000000000000", 20596 => "0000000000000000", 20597 => "0000000000000000", 20598 => "0000000000000000", 20599 => "0000000000000000", 20600 => "0000000000000000", 20601 => "0000000000000000", 20602 => "0000000000000000", 20603 => "0000000000000000", 20604 => "0000000000000000", 20605 => "0000000000000000", 20606 => "0000000000000000", 20607 => "0000000000000000", 20608 => "0000000000000000", 20609 => "0000000000000000", 20610 => "0000000000000000", 20611 => "0000000000000000", 20612 => "0000000000000000", 20613 => "0000000000000000", 20614 => "0000000000000000", 20615 => "0000000000000000", 20616 => "0000000000000000", 20617 => "0000000000000000", 20618 => "0000000000000000", 20619 => "0000000000000000", 20620 => "0000000000000000", 20621 => "0000000000000000", 20622 => "0000000000000000", 20623 => "0000000000000000", 20624 => "0000000000000000", 20625 => "0000000000000000", 20626 => "0000000000000000", 20627 => "0000000000000000", 20628 => "0000000000000000", 20629 => "0000000000000000", 20630 => "0000000000000000", 20631 => "0000000000000000", 20632 => "0000000000000000", 20633 => "0000000000000000", 20634 => "0000000000000000", 20635 => "0000000000000000", 20636 => "0000000000000000", 20637 => "0000000000000000", 20638 => "0000000000000000", 20639 => "0000000000000000", 20640 => "0000000000000000", 20641 => "0000000000000000", 20642 => "0000000000000000", 20643 => "0000000000000000", 20644 => "0000000000000000", 20645 => "0000000000000000", 20646 => "0000000000000000", 20647 => "0000000000000000", 20648 => "0000000000000000", 20649 => "0000000000000000", 20650 => "0000000000000000", 20651 => "0000000000000000", 20652 => "0000000000000000", 20653 => "0000000000000000", 20654 => "0000000000000000", 20655 => "0000000000000000", 20656 => "0000000000000000", 20657 => "0000000000000000", 20658 => "0000000000000000", 20659 => "0000000000000000", 20660 => "0000000000000000", 20661 => "0000000000000000", 20662 => "0000000000000000", 20663 => "0000000000000000", 20664 => "0000000000000000", 20665 => "0000000000000000", 20666 => "0000000000000000", 20667 => "0000000000000000", 20668 => "0000000000000000", 20669 => "0000000000000000", 20670 => "0000000000000000", 20671 => "0000000000000000", 20672 => "0000000000000000", 20673 => "0000000000000000", 20674 => "0000000000000000", 20675 => "0000000000000000", 20676 => "0000000000000000", 20677 => "0000000000000000", 20678 => "0000000000000000", 20679 => "0000000000000000", 20680 => "0000000000000000", 20681 => "0000000000000000", 20682 => "0000000000000000", 20683 => "0000000000000000", 20684 => "0000000000000000", 20685 => "0000000000000000", 20686 => "0000000000000000", 20687 => "0000000000000000", 20688 => "0000000000000000", 20689 => "0000000000000000", 20690 => "0000000000000000", 20691 => "0000000000000000", 20692 => "0000000000000000", 20693 => "0000000000000000", 20694 => "0000000000000000", 20695 => "0000000000000000", 20696 => "0000000000000000", 20697 => "0000000000000000", 20698 => "0000000000000000", 20699 => "0000000000000000", 20700 => "0000000000000000", 20701 => "0000000000000000", 20702 => "0000000000000000", 20703 => "0000000000000000", 20704 => "0000000000000000", 20705 => "0000000000000000", 20706 => "0000000000000000", 20707 => "0000000000000000", 20708 => "0000000000000000", 20709 => "0000000000000000", 20710 => "0000000000000000", 20711 => "0000000000000000", 20712 => "0000000000000000", 20713 => "0000000000000000", 20714 => "0000000000000000", 20715 => "0000000000000000", 20716 => "0000000000000000", 20717 => "0000000000000000", 20718 => "0000000000000000", 20719 => "0000000000000000", 20720 => "0000000000000000", 20721 => "0000000000000000", 20722 => "0000000000000000", 20723 => "0000000000000000", 20724 => "0000000000000000", 20725 => "0000000000000000", 20726 => "0000000000000000", 20727 => "0000000000000000", 20728 => "0000000000000000", 20729 => "0000000000000000", 20730 => "0000000000000000", 20731 => "0000000000000000", 20732 => "0000000000000000", 20733 => "0000000000000000", 20734 => "0000000000000000", 20735 => "0000000000000000", 20736 => "0000000000000000", 20737 => "0000000000000000", 20738 => "0000000000000000", 20739 => "0000000000000000", 20740 => "0000000000000000", 20741 => "0000000000000000", 20742 => "0000000000000000", 20743 => "0000000000000000", 20744 => "0000000000000000", 20745 => "0000000000000000", 20746 => "0000000000000000", 20747 => "0000000000000000", 20748 => "0000000000000000", 20749 => "0000000000000000", 20750 => "0000000000000000", 20751 => "0000000000000000", 20752 => "0000000000000000", 20753 => "0000000000000000", 20754 => "0000000000000000", 20755 => "0000000000000000", 20756 => "0000000000000000", 20757 => "0000000000000000", 20758 => "0000000000000000", 20759 => "0000000000000000", 20760 => "0000000000000000", 20761 => "0000000000000000", 20762 => "0000000000000000", 20763 => "0000000000000000", 20764 => "0000000000000000", 20765 => "0000000000000000", 20766 => "0000000000000000", 20767 => "0000000000000000", 20768 => "0000000000000000", 20769 => "0000000000000000", 20770 => "0000000000000000", 20771 => "0000000000000000", 20772 => "0000000000000000", 20773 => "0000000000000000", 20774 => "0000000000000000", 20775 => "0000000000000000", 20776 => "0000000000000000", 20777 => "0000000000000000", 20778 => "0000000000000000", 20779 => "0000000000000000", 20780 => "0000000000000000", 20781 => "0000000000000000", 20782 => "0000000000000000", 20783 => "0000000000000000", 20784 => "0000000000000000", 20785 => "0000000000000000", 20786 => "0000000000000000", 20787 => "0000000000000000", 20788 => "0000000000000000", 20789 => "0000000000000000", 20790 => "0000000000000000", 20791 => "0000000000000000", 20792 => "0000000000000000", 20793 => "0000000000000000", 20794 => "0000000000000000", 20795 => "0000000000000000", 20796 => "0000000000000000", 20797 => "0000000000000000", 20798 => "0000000000000000", 20799 => "0000000000000000", 20800 => "0000000000000000", 20801 => "0000000000000000", 20802 => "0000000000000000", 20803 => "0000000000000000", 20804 => "0000000000000000", 20805 => "0000000000000000", 20806 => "0000000000000000", 20807 => "0000000000000000", 20808 => "0000000000000000", 20809 => "0000000000000000", 20810 => "0000000000000000", 20811 => "0000000000000000", 20812 => "0000000000000000", 20813 => "0000000000000000", 20814 => "0000000000000000", 20815 => "0000000000000000", 20816 => "0000000000000000", 20817 => "0000000000000000", 20818 => "0000000000000000", 20819 => "0000000000000000", 20820 => "0000000000000000", 20821 => "0000000000000000", 20822 => "0000000000000000", 20823 => "0000000000000000", 20824 => "0000000000000000", 20825 => "0000000000000000", 20826 => "0000000000000000", 20827 => "0000000000000000", 20828 => "0000000000000000", 20829 => "0000000000000000", 20830 => "0000000000000000", 20831 => "0000000000000000", 20832 => "0000000000000000", 20833 => "0000000000000000", 20834 => "0000000000000000", 20835 => "0000000000000000", 20836 => "0000000000000000", 20837 => "0000000000000000", 20838 => "0000000000000000", 20839 => "0000000000000000", 20840 => "0000000000000000", 20841 => "0000000000000000", 20842 => "0000000000000000", 20843 => "0000000000000000", 20844 => "0000000000000000", 20845 => "0000000000000000", 20846 => "0000000000000000", 20847 => "0000000000000000", 20848 => "0000000000000000", 20849 => "0000000000000000", 20850 => "0000000000000000", 20851 => "0000000000000000", 20852 => "0000000000000000", 20853 => "0000000000000000", 20854 => "0000000000000000", 20855 => "0000000000000000", 20856 => "0000000000000000", 20857 => "0000000000000000", 20858 => "0000000000000000", 20859 => "0000000000000000", 20860 => "0000000000000000", 20861 => "0000000000000000", 20862 => "0000000000000000", 20863 => "0000000000000000", 20864 => "0000000000000000", 20865 => "0000000000000000", 20866 => "0000000000000000", 20867 => "0000000000000000", 20868 => "0000000000000000", 20869 => "0000000000000000", 20870 => "0000000000000000", 20871 => "0000000000000000", 20872 => "0000000000000000", 20873 => "0000000000000000", 20874 => "0000000000000000", 20875 => "0000000000000000", 20876 => "0000000000000000", 20877 => "0000000000000000", 20878 => "0000000000000000", 20879 => "0000000000000000", 20880 => "0000000000000000", 20881 => "0000000000000000", 20882 => "0000000000000000", 20883 => "0000000000000000", 20884 => "0000000000000000", 20885 => "0000000000000000", 20886 => "0000000000000000", 20887 => "0000000000000000", 20888 => "0000000000000000", 20889 => "0000000000000000", 20890 => "0000000000000000", 20891 => "0000000000000000", 20892 => "0000000000000000", 20893 => "0000000000000000", 20894 => "0000000000000000", 20895 => "0000000000000000", 20896 => "0000000000000000", 20897 => "0000000000000000", 20898 => "0000000000000000", 20899 => "0000000000000000", 20900 => "0000000000000000", 20901 => "0000000000000000", 20902 => "0000000000000000", 20903 => "0000000000000000", 20904 => "0000000000000000", 20905 => "0000000000000000", 20906 => "0000000000000000", 20907 => "0000000000000000", 20908 => "0000000000000000", 20909 => "0000000000000000", 20910 => "0000000000000000", 20911 => "0000000000000000", 20912 => "0000000000000000", 20913 => "0000000000000000", 20914 => "0000000000000000", 20915 => "0000000000000000", 20916 => "0000000000000000", 20917 => "0000000000000000", 20918 => "0000000000000000", 20919 => "0000000000000000", 20920 => "0000000000000000", 20921 => "0000000000000000", 20922 => "0000000000000000", 20923 => "0000000000000000", 20924 => "0000000000000000", 20925 => "0000000000000000", 20926 => "0000000000000000", 20927 => "0000000000000000", 20928 => "0000000000000000", 20929 => "0000000000000000", 20930 => "0000000000000000", 20931 => "0000000000000000", 20932 => "0000000000000000", 20933 => "0000000000000000", 20934 => "0000000000000000", 20935 => "0000000000000000", 20936 => "0000000000000000", 20937 => "0000000000000000", 20938 => "0000000000000000", 20939 => "0000000000000000", 20940 => "0000000000000000", 20941 => "0000000000000000", 20942 => "0000000000000000", 20943 => "0000000000000000", 20944 => "0000000000000000", 20945 => "0000000000000000", 20946 => "0000000000000000", 20947 => "0000000000000000", 20948 => "0000000000000000", 20949 => "0000000000000000", 20950 => "0000000000000000", 20951 => "0000000000000000", 20952 => "0000000000000000", 20953 => "0000000000000000", 20954 => "0000000000000000", 20955 => "0000000000000000", 20956 => "0000000000000000", 20957 => "0000000000000000", 20958 => "0000000000000000", 20959 => "0000000000000000", 20960 => "0000000000000000", 20961 => "0000000000000000", 20962 => "0000000000000000", 20963 => "0000000000000000", 20964 => "0000000000000000", 20965 => "0000000000000000", 20966 => "0000000000000000", 20967 => "0000000000000000", 20968 => "0000000000000000", 20969 => "0000000000000000", 20970 => "0000000000000000", 20971 => "0000000000000000", 20972 => "0000000000000000", 20973 => "0000000000000000", 20974 => "0000000000000000", 20975 => "0000000000000000", 20976 => "0000000000000000", 20977 => "0000000000000000", 20978 => "0000000000000000", 20979 => "0000000000000000", 20980 => "0000000000000000", 20981 => "0000000000000000", 20982 => "0000000000000000", 20983 => "0000000000000000", 20984 => "0000000000000000", 20985 => "0000000000000000", 20986 => "0000000000000000", 20987 => "0000000000000000", 20988 => "0000000000000000", 20989 => "0000000000000000", 20990 => "0000000000000000", 20991 => "0000000000000000", 20992 => "0000000000000000", 20993 => "0000000000000000", 20994 => "0000000000000000", 20995 => "0000000000000000", 20996 => "0000000000000000", 20997 => "0000000000000000", 20998 => "0000000000000000", 20999 => "0000000000000000", 21000 => "0000000000000000", 21001 => "0000000000000000", 21002 => "0000000000000000", 21003 => "0000000000000000", 21004 => "0000000000000000", 21005 => "0000000000000000", 21006 => "0000000000000000", 21007 => "0000000000000000", 21008 => "0000000000000000", 21009 => "0000000000000000", 21010 => "0000000000000000", 21011 => "0000000000000000", 21012 => "0000000000000000", 21013 => "0000000000000000", 21014 => "0000000000000000", 21015 => "0000000000000000", 21016 => "0000000000000000", 21017 => "0000000000000000", 21018 => "0000000000000000", 21019 => "0000000000000000", 21020 => "0000000000000000", 21021 => "0000000000000000", 21022 => "0000000000000000", 21023 => "0000000000000000", 21024 => "0000000000000000", 21025 => "0000000000000000", 21026 => "0000000000000000", 21027 => "0000000000000000", 21028 => "0000000000000000", 21029 => "0000000000000000", 21030 => "0000000000000000", 21031 => "0000000000000000", 21032 => "0000000000000000", 21033 => "0000000000000000", 21034 => "0000000000000000", 21035 => "0000000000000000", 21036 => "0000000000000000", 21037 => "0000000000000000", 21038 => "0000000000000000", 21039 => "0000000000000000", 21040 => "0000000000000000", 21041 => "0000000000000000", 21042 => "0000000000000000", 21043 => "0000000000000000", 21044 => "0000000000000000", 21045 => "0000000000000000", 21046 => "0000000000000000", 21047 => "0000000000000000", 21048 => "0000000000000000", 21049 => "0000000000000000", 21050 => "0000000000000000", 21051 => "0000000000000000", 21052 => "0000000000000000", 21053 => "0000000000000000", 21054 => "0000000000000000", 21055 => "0000000000000000", 21056 => "0000000000000000", 21057 => "0000000000000000", 21058 => "0000000000000000", 21059 => "0000000000000000", 21060 => "0000000000000000", 21061 => "0000000000000000", 21062 => "0000000000000000", 21063 => "0000000000000000", 21064 => "0000000000000000", 21065 => "0000000000000000", 21066 => "0000000000000000", 21067 => "0000000000000000", 21068 => "0000000000000000", 21069 => "0000000000000000", 21070 => "0000000000000000", 21071 => "0000000000000000", 21072 => "0000000000000000", 21073 => "0000000000000000", 21074 => "0000000000000000", 21075 => "0000000000000000", 21076 => "0000000000000000", 21077 => "0000000000000000", 21078 => "0000000000000000", 21079 => "0000000000000000", 21080 => "0000000000000000", 21081 => "0000000000000000", 21082 => "0000000000000000", 21083 => "0000000000000000", 21084 => "0000000000000000", 21085 => "0000000000000000", 21086 => "0000000000000000", 21087 => "0000000000000000", 21088 => "0000000000000000", 21089 => "0000000000000000", 21090 => "0000000000000000", 21091 => "0000000000000000", 21092 => "0000000000000000", 21093 => "0000000000000000", 21094 => "0000000000000000", 21095 => "0000000000000000", 21096 => "0000000000000000", 21097 => "0000000000000000", 21098 => "0000000000000000", 21099 => "0000000000000000", 21100 => "0000000000000000", 21101 => "0000000000000000", 21102 => "0000000000000000", 21103 => "0000000000000000", 21104 => "0000000000000000", 21105 => "0000000000000000", 21106 => "0000000000000000", 21107 => "0000000000000000", 21108 => "0000000000000000", 21109 => "0000000000000000", 21110 => "0000000000000000", 21111 => "0000000000000000", 21112 => "0000000000000000", 21113 => "0000000000000000", 21114 => "0000000000000000", 21115 => "0000000000000000", 21116 => "0000000000000000", 21117 => "0000000000000000", 21118 => "0000000000000000", 21119 => "0000000000000000", 21120 => "0000000000000000", 21121 => "0000000000000000", 21122 => "0000000000000000", 21123 => "0000000000000000", 21124 => "0000000000000000", 21125 => "0000000000000000", 21126 => "0000000000000000", 21127 => "0000000000000000", 21128 => "0000000000000000", 21129 => "0000000000000000", 21130 => "0000000000000000", 21131 => "0000000000000000", 21132 => "0000000000000000", 21133 => "0000000000000000", 21134 => "0000000000000000", 21135 => "0000000000000000", 21136 => "0000000000000000", 21137 => "0000000000000000", 21138 => "0000000000000000", 21139 => "0000000000000000", 21140 => "0000000000000000", 21141 => "0000000000000000", 21142 => "0000000000000000", 21143 => "0000000000000000", 21144 => "0000000000000000", 21145 => "0000000000000000", 21146 => "0000000000000000", 21147 => "0000000000000000", 21148 => "0000000000000000", 21149 => "0000000000000000", 21150 => "0000000000000000", 21151 => "0000000000000000", 21152 => "0000000000000000", 21153 => "0000000000000000", 21154 => "0000000000000000", 21155 => "0000000000000000", 21156 => "0000000000000000", 21157 => "0000000000000000", 21158 => "0000000000000000", 21159 => "0000000000000000", 21160 => "0000000000000000", 21161 => "0000000000000000", 21162 => "0000000000000000", 21163 => "0000000000000000", 21164 => "0000000000000000", 21165 => "0000000000000000", 21166 => "0000000000000000", 21167 => "0000000000000000", 21168 => "0000000000000000", 21169 => "0000000000000000", 21170 => "0000000000000000", 21171 => "0000000000000000", 21172 => "0000000000000000", 21173 => "0000000000000000", 21174 => "0000000000000000", 21175 => "0000000000000000", 21176 => "0000000000000000", 21177 => "0000000000000000", 21178 => "0000000000000000", 21179 => "0000000000000000", 21180 => "0000000000000000", 21181 => "0000000000000000", 21182 => "0000000000000000", 21183 => "0000000000000000", 21184 => "0000000000000000", 21185 => "0000000000000000", 21186 => "0000000000000000", 21187 => "0000000000000000", 21188 => "0000000000000000", 21189 => "0000000000000000", 21190 => "0000000000000000", 21191 => "0000000000000000", 21192 => "0000000000000000", 21193 => "0000000000000000", 21194 => "0000000000000000", 21195 => "0000000000000000", 21196 => "0000000000000000", 21197 => "0000000000000000", 21198 => "0000000000000000", 21199 => "0000000000000000", 21200 => "0000000000000000", 21201 => "0000000000000000", 21202 => "0000000000000000", 21203 => "0000000000000000", 21204 => "0000000000000000", 21205 => "0000000000000000", 21206 => "0000000000000000", 21207 => "0000000000000000", 21208 => "0000000000000000", 21209 => "0000000000000000", 21210 => "0000000000000000", 21211 => "0000000000000000", 21212 => "0000000000000000", 21213 => "0000000000000000", 21214 => "0000000000000000", 21215 => "0000000000000000", 21216 => "0000000000000000", 21217 => "0000000000000000", 21218 => "0000000000000000", 21219 => "0000000000000000", 21220 => "0000000000000000", 21221 => "0000000000000000", 21222 => "0000000000000000", 21223 => "0000000000000000", 21224 => "0000000000000000", 21225 => "0000000000000000", 21226 => "0000000000000000", 21227 => "0000000000000000", 21228 => "0000000000000000", 21229 => "0000000000000000", 21230 => "0000000000000000", 21231 => "0000000000000000", 21232 => "0000000000000000", 21233 => "0000000000000000", 21234 => "0000000000000000", 21235 => "0000000000000000", 21236 => "0000000000000000", 21237 => "0000000000000000", 21238 => "0000000000000000", 21239 => "0000000000000000", 21240 => "0000000000000000", 21241 => "0000000000000000", 21242 => "0000000000000000", 21243 => "0000000000000000", 21244 => "0000000000000000", 21245 => "0000000000000000", 21246 => "0000000000000000", 21247 => "0000000000000000", 21248 => "0000000000000000", 21249 => "0000000000000000", 21250 => "0000000000000000", 21251 => "0000000000000000", 21252 => "0000000000000000", 21253 => "0000000000000000", 21254 => "0000000000000000", 21255 => "0000000000000000", 21256 => "0000000000000000", 21257 => "0000000000000000", 21258 => "0000000000000000", 21259 => "0000000000000000", 21260 => "0000000000000000", 21261 => "0000000000000000", 21262 => "0000000000000000", 21263 => "0000000000000000", 21264 => "0000000000000000", 21265 => "0000000000000000", 21266 => "0000000000000000", 21267 => "0000000000000000", 21268 => "0000000000000000", 21269 => "0000000000000000", 21270 => "0000000000000000", 21271 => "0000000000000000", 21272 => "0000000000000000", 21273 => "0000000000000000", 21274 => "0000000000000000", 21275 => "0000000000000000", 21276 => "0000000000000000", 21277 => "0000000000000000", 21278 => "0000000000000000", 21279 => "0000000000000000", 21280 => "0000000000000000", 21281 => "0000000000000000", 21282 => "0000000000000000", 21283 => "0000000000000000", 21284 => "0000000000000000", 21285 => "0000000000000000", 21286 => "0000000000000000", 21287 => "0000000000000000", 21288 => "0000000000000000", 21289 => "0000000000000000", 21290 => "0000000000000000", 21291 => "0000000000000000", 21292 => "0000000000000000", 21293 => "0000000000000000", 21294 => "0000000000000000", 21295 => "0000000000000000", 21296 => "0000000000000000", 21297 => "0000000000000000", 21298 => "0000000000000000", 21299 => "0000000000000000", 21300 => "0000000000000000", 21301 => "0000000000000000", 21302 => "0000000000000000", 21303 => "0000000000000000", 21304 => "0000000000000000", 21305 => "0000000000000000", 21306 => "0000000000000000", 21307 => "0000000000000000", 21308 => "0000000000000000", 21309 => "0000000000000000", 21310 => "0000000000000000", 21311 => "0000000000000000", 21312 => "0000000000000000", 21313 => "0000000000000000", 21314 => "0000000000000000", 21315 => "0000000000000000", 21316 => "0000000000000000", 21317 => "0000000000000000", 21318 => "0000000000000000", 21319 => "0000000000000000", 21320 => "0000000000000000", 21321 => "0000000000000000", 21322 => "0000000000000000", 21323 => "0000000000000000", 21324 => "0000000000000000", 21325 => "0000000000000000", 21326 => "0000000000000000", 21327 => "0000000000000000", 21328 => "0000000000000000", 21329 => "0000000000000000", 21330 => "0000000000000000", 21331 => "0000000000000000", 21332 => "0000000000000000", 21333 => "0000000000000000", 21334 => "0000000000000000", 21335 => "0000000000000000", 21336 => "0000000000000000", 21337 => "0000000000000000", 21338 => "0000000000000000", 21339 => "0000000000000000", 21340 => "0000000000000000", 21341 => "0000000000000000", 21342 => "0000000000000000", 21343 => "0000000000000000", 21344 => "0000000000000000", 21345 => "0000000000000000", 21346 => "0000000000000000", 21347 => "0000000000000000", 21348 => "0000000000000000", 21349 => "0000000000000000", 21350 => "0000000000000000", 21351 => "0000000000000000", 21352 => "0000000000000000", 21353 => "0000000000000000", 21354 => "0000000000000000", 21355 => "0000000000000000", 21356 => "0000000000000000", 21357 => "0000000000000000", 21358 => "0000000000000000", 21359 => "0000000000000000", 21360 => "0000000000000000", 21361 => "0000000000000000", 21362 => "0000000000000000", 21363 => "0000000000000000", 21364 => "0000000000000000", 21365 => "0000000000000000", 21366 => "0000000000000000", 21367 => "0000000000000000", 21368 => "0000000000000000", 21369 => "0000000000000000", 21370 => "0000000000000000", 21371 => "0000000000000000", 21372 => "0000000000000000", 21373 => "0000000000000000", 21374 => "0000000000000000", 21375 => "0000000000000000", 21376 => "0000000000000000", 21377 => "0000000000000000", 21378 => "0000000000000000", 21379 => "0000000000000000", 21380 => "0000000000000000", 21381 => "0000000000000000", 21382 => "0000000000000000", 21383 => "0000000000000000", 21384 => "0000000000000000", 21385 => "0000000000000000", 21386 => "0000000000000000", 21387 => "0000000000000000", 21388 => "0000000000000000", 21389 => "0000000000000000", 21390 => "0000000000000000", 21391 => "0000000000000000", 21392 => "0000000000000000", 21393 => "0000000000000000", 21394 => "0000000000000000", 21395 => "0000000000000000", 21396 => "0000000000000000", 21397 => "0000000000000000", 21398 => "0000000000000000", 21399 => "0000000000000000", 21400 => "0000000000000000", 21401 => "0000000000000000", 21402 => "0000000000000000", 21403 => "0000000000000000", 21404 => "0000000000000000", 21405 => "0000000000000000", 21406 => "0000000000000000", 21407 => "0000000000000000", 21408 => "0000000000000000", 21409 => "0000000000000000", 21410 => "0000000000000000", 21411 => "0000000000000000", 21412 => "0000000000000000", 21413 => "0000000000000000", 21414 => "0000000000000000", 21415 => "0000000000000000", 21416 => "0000000000000000", 21417 => "0000000000000000", 21418 => "0000000000000000", 21419 => "0000000000000000", 21420 => "0000000000000000", 21421 => "0000000000000000", 21422 => "0000000000000000", 21423 => "0000000000000000", 21424 => "0000000000000000", 21425 => "0000000000000000", 21426 => "0000000000000000", 21427 => "0000000000000000", 21428 => "0000000000000000", 21429 => "0000000000000000", 21430 => "0000000000000000", 21431 => "0000000000000000", 21432 => "0000000000000000", 21433 => "0000000000000000", 21434 => "0000000000000000", 21435 => "0000000000000000", 21436 => "0000000000000000", 21437 => "0000000000000000", 21438 => "0000000000000000", 21439 => "0000000000000000", 21440 => "0000000000000000", 21441 => "0000000000000000", 21442 => "0000000000000000", 21443 => "0000000000000000", 21444 => "0000000000000000", 21445 => "0000000000000000", 21446 => "0000000000000000", 21447 => "0000000000000000", 21448 => "0000000000000000", 21449 => "0000000000000000", 21450 => "0000000000000000", 21451 => "0000000000000000", 21452 => "0000000000000000", 21453 => "0000000000000000", 21454 => "0000000000000000", 21455 => "0000000000000000", 21456 => "0000000000000000", 21457 => "0000000000000000", 21458 => "0000000000000000", 21459 => "0000000000000000", 21460 => "0000000000000000", 21461 => "0000000000000000", 21462 => "0000000000000000", 21463 => "0000000000000000", 21464 => "0000000000000000", 21465 => "0000000000000000", 21466 => "0000000000000000", 21467 => "0000000000000000", 21468 => "0000000000000000", 21469 => "0000000000000000", 21470 => "0000000000000000", 21471 => "0000000000000000", 21472 => "0000000000000000", 21473 => "0000000000000000", 21474 => "0000000000000000", 21475 => "0000000000000000", 21476 => "0000000000000000", 21477 => "0000000000000000", 21478 => "0000000000000000", 21479 => "0000000000000000", 21480 => "0000000000000000", 21481 => "0000000000000000", 21482 => "0000000000000000", 21483 => "0000000000000000", 21484 => "0000000000000000", 21485 => "0000000000000000", 21486 => "0000000000000000", 21487 => "0000000000000000", 21488 => "0000000000000000", 21489 => "0000000000000000", 21490 => "0000000000000000", 21491 => "0000000000000000", 21492 => "0000000000000000", 21493 => "0000000000000000", 21494 => "0000000000000000", 21495 => "0000000000000000", 21496 => "0000000000000000", 21497 => "0000000000000000", 21498 => "0000000000000000", 21499 => "0000000000000000", 21500 => "0000000000000000", 21501 => "0000000000000000", 21502 => "0000000000000000", 21503 => "0000000000000000", 21504 => "0000000000000000", 21505 => "0000000000000000", 21506 => "0000000000000000", 21507 => "0000000000000000", 21508 => "0000000000000000", 21509 => "0000000000000000", 21510 => "0000000000000000", 21511 => "0000000000000000", 21512 => "0000000000000000", 21513 => "0000000000000000", 21514 => "0000000000000000", 21515 => "0000000000000000", 21516 => "0000000000000000", 21517 => "0000000000000000", 21518 => "0000000000000000", 21519 => "0000000000000000", 21520 => "0000000000000000", 21521 => "0000000000000000", 21522 => "0000000000000000", 21523 => "0000000000000000", 21524 => "0000000000000000", 21525 => "0000000000000000", 21526 => "0000000000000000", 21527 => "0000000000000000", 21528 => "0000000000000000", 21529 => "0000000000000000", 21530 => "0000000000000000", 21531 => "0000000000000000", 21532 => "0000000000000000", 21533 => "0000000000000000", 21534 => "0000000000000000", 21535 => "0000000000000000", 21536 => "0000000000000000", 21537 => "0000000000000000", 21538 => "0000000000000000", 21539 => "0000000000000000", 21540 => "0000000000000000", 21541 => "0000000000000000", 21542 => "0000000000000000", 21543 => "0000000000000000", 21544 => "0000000000000000", 21545 => "0000000000000000", 21546 => "0000000000000000", 21547 => "0000000000000000", 21548 => "0000000000000000", 21549 => "0000000000000000", 21550 => "0000000000000000", 21551 => "0000000000000000", 21552 => "0000000000000000", 21553 => "0000000000000000", 21554 => "0000000000000000", 21555 => "0000000000000000", 21556 => "0000000000000000", 21557 => "0000000000000000", 21558 => "0000000000000000", 21559 => "0000000000000000", 21560 => "0000000000000000", 21561 => "0000000000000000", 21562 => "0000000000000000", 21563 => "0000000000000000", 21564 => "0000000000000000", 21565 => "0000000000000000", 21566 => "0000000000000000", 21567 => "0000000000000000", 21568 => "0000000000000000", 21569 => "0000000000000000", 21570 => "0000000000000000", 21571 => "0000000000000000", 21572 => "0000000000000000", 21573 => "0000000000000000", 21574 => "0000000000000000", 21575 => "0000000000000000", 21576 => "0000000000000000", 21577 => "0000000000000000", 21578 => "0000000000000000", 21579 => "0000000000000000", 21580 => "0000000000000000", 21581 => "0000000000000000", 21582 => "0000000000000000", 21583 => "0000000000000000", 21584 => "0000000000000000", 21585 => "0000000000000000", 21586 => "0000000000000000", 21587 => "0000000000000000", 21588 => "0000000000000000", 21589 => "0000000000000000", 21590 => "0000000000000000", 21591 => "0000000000000000", 21592 => "0000000000000000", 21593 => "0000000000000000", 21594 => "0000000000000000", 21595 => "0000000000000000", 21596 => "0000000000000000", 21597 => "0000000000000000", 21598 => "0000000000000000", 21599 => "0000000000000000", 21600 => "0000000000000000", 21601 => "0000000000000000", 21602 => "0000000000000000", 21603 => "0000000000000000", 21604 => "0000000000000000", 21605 => "0000000000000000", 21606 => "0000000000000000", 21607 => "0000000000000000", 21608 => "0000000000000000", 21609 => "0000000000000000", 21610 => "0000000000000000", 21611 => "0000000000000000", 21612 => "0000000000000000", 21613 => "0000000000000000", 21614 => "0000000000000000", 21615 => "0000000000000000", 21616 => "0000000000000000", 21617 => "0000000000000000", 21618 => "0000000000000000", 21619 => "0000000000000000", 21620 => "0000000000000000", 21621 => "0000000000000000", 21622 => "0000000000000000", 21623 => "0000000000000000", 21624 => "0000000000000000", 21625 => "0000000000000000", 21626 => "0000000000000000", 21627 => "0000000000000000", 21628 => "0000000000000000", 21629 => "0000000000000000", 21630 => "0000000000000000", 21631 => "0000000000000000", 21632 => "0000000000000000", 21633 => "0000000000000000", 21634 => "0000000000000000", 21635 => "0000000000000000", 21636 => "0000000000000000", 21637 => "0000000000000000", 21638 => "0000000000000000", 21639 => "0000000000000000", 21640 => "0000000000000000", 21641 => "0000000000000000", 21642 => "0000000000000000", 21643 => "0000000000000000", 21644 => "0000000000000000", 21645 => "0000000000000000", 21646 => "0000000000000000", 21647 => "0000000000000000", 21648 => "0000000000000000", 21649 => "0000000000000000", 21650 => "0000000000000000", 21651 => "0000000000000000", 21652 => "0000000000000000", 21653 => "0000000000000000", 21654 => "0000000000000000", 21655 => "0000000000000000", 21656 => "0000000000000000", 21657 => "0000000000000000", 21658 => "0000000000000000", 21659 => "0000000000000000", 21660 => "0000000000000000", 21661 => "0000000000000000", 21662 => "0000000000000000", 21663 => "0000000000000000", 21664 => "0000000000000000", 21665 => "0000000000000000", 21666 => "0000000000000000", 21667 => "0000000000000000", 21668 => "0000000000000000", 21669 => "0000000000000000", 21670 => "0000000000000000", 21671 => "0000000000000000", 21672 => "0000000000000000", 21673 => "0000000000000000", 21674 => "0000000000000000", 21675 => "0000000000000000", 21676 => "0000000000000000", 21677 => "0000000000000000", 21678 => "0000000000000000", 21679 => "0000000000000000", 21680 => "0000000000000000", 21681 => "0000000000000000", 21682 => "0000000000000000", 21683 => "0000000000000000", 21684 => "0000000000000000", 21685 => "0000000000000000", 21686 => "0000000000000000", 21687 => "0000000000000000", 21688 => "0000000000000000", 21689 => "0000000000000000", 21690 => "0000000000000000", 21691 => "0000000000000000", 21692 => "0000000000000000", 21693 => "0000000000000000", 21694 => "0000000000000000", 21695 => "0000000000000000", 21696 => "0000000000000000", 21697 => "0000000000000000", 21698 => "0000000000000000", 21699 => "0000000000000000", 21700 => "0000000000000000", 21701 => "0000000000000000", 21702 => "0000000000000000", 21703 => "0000000000000000", 21704 => "0000000000000000", 21705 => "0000000000000000", 21706 => "0000000000000000", 21707 => "0000000000000000", 21708 => "0000000000000000", 21709 => "0000000000000000", 21710 => "0000000000000000", 21711 => "0000000000000000", 21712 => "0000000000000000", 21713 => "0000000000000000", 21714 => "0000000000000000", 21715 => "0000000000000000", 21716 => "0000000000000000", 21717 => "0000000000000000", 21718 => "0000000000000000", 21719 => "0000000000000000", 21720 => "0000000000000000", 21721 => "0000000000000000", 21722 => "0000000000000000", 21723 => "0000000000000000", 21724 => "0000000000000000", 21725 => "0000000000000000", 21726 => "0000000000000000", 21727 => "0000000000000000", 21728 => "0000000000000000", 21729 => "0000000000000000", 21730 => "0000000000000000", 21731 => "0000000000000000", 21732 => "0000000000000000", 21733 => "0000000000000000", 21734 => "0000000000000000", 21735 => "0000000000000000", 21736 => "0000000000000000", 21737 => "0000000000000000", 21738 => "0000000000000000", 21739 => "0000000000000000", 21740 => "0000000000000000", 21741 => "0000000000000000", 21742 => "0000000000000000", 21743 => "0000000000000000", 21744 => "0000000000000000", 21745 => "0000000000000000", 21746 => "0000000000000000", 21747 => "0000000000000000", 21748 => "0000000000000000", 21749 => "0000000000000000", 21750 => "0000000000000000", 21751 => "0000000000000000", 21752 => "0000000000000000", 21753 => "0000000000000000", 21754 => "0000000000000000", 21755 => "0000000000000000", 21756 => "0000000000000000", 21757 => "0000000000000000", 21758 => "0000000000000000", 21759 => "0000000000000000", 21760 => "0000000000000000", 21761 => "0000000000000000", 21762 => "0000000000000000", 21763 => "0000000000000000", 21764 => "0000000000000000", 21765 => "0000000000000000", 21766 => "0000000000000000", 21767 => "0000000000000000", 21768 => "0000000000000000", 21769 => "0000000000000000", 21770 => "0000000000000000", 21771 => "0000000000000000", 21772 => "0000000000000000", 21773 => "0000000000000000", 21774 => "0000000000000000", 21775 => "0000000000000000", 21776 => "0000000000000000", 21777 => "0000000000000000", 21778 => "0000000000000000", 21779 => "0000000000000000", 21780 => "0000000000000000", 21781 => "0000000000000000", 21782 => "0000000000000000", 21783 => "0000000000000000", 21784 => "0000000000000000", 21785 => "0000000000000000", 21786 => "0000000000000000", 21787 => "0000000000000000", 21788 => "0000000000000000", 21789 => "0000000000000000", 21790 => "0000000000000000", 21791 => "0000000000000000", 21792 => "0000000000000000", 21793 => "0000000000000000", 21794 => "0000000000000000", 21795 => "0000000000000000", 21796 => "0000000000000000", 21797 => "0000000000000000", 21798 => "0000000000000000", 21799 => "0000000000000000", 21800 => "0000000000000000", 21801 => "0000000000000000", 21802 => "0000000000000000", 21803 => "0000000000000000", 21804 => "0000000000000000", 21805 => "0000000000000000", 21806 => "0000000000000000", 21807 => "0000000000000000", 21808 => "0000000000000000", 21809 => "0000000000000000", 21810 => "0000000000000000", 21811 => "0000000000000000", 21812 => "0000000000000000", 21813 => "0000000000000000", 21814 => "0000000000000000", 21815 => "0000000000000000", 21816 => "0000000000000000", 21817 => "0000000000000000", 21818 => "0000000000000000", 21819 => "0000000000000000", 21820 => "0000000000000000", 21821 => "0000000000000000", 21822 => "0000000000000000", 21823 => "0000000000000000", 21824 => "0000000000000000", 21825 => "0000000000000000", 21826 => "0000000000000000", 21827 => "0000000000000000", 21828 => "0000000000000000", 21829 => "0000000000000000", 21830 => "0000000000000000", 21831 => "0000000000000000", 21832 => "0000000000000000", 21833 => "0000000000000000", 21834 => "0000000000000000", 21835 => "0000000000000000", 21836 => "0000000000000000", 21837 => "0000000000000000", 21838 => "0000000000000000", 21839 => "0000000000000000", 21840 => "0000000000000000", 21841 => "0000000000000000", 21842 => "0000000000000000", 21843 => "0000000000000000", 21844 => "0000000000000000", 21845 => "0000000000000000", 21846 => "0000000000000000", 21847 => "0000000000000000", 21848 => "0000000000000000", 21849 => "0000000000000000", 21850 => "0000000000000000", 21851 => "0000000000000000", 21852 => "0000000000000000", 21853 => "0000000000000000", 21854 => "0000000000000000", 21855 => "0000000000000000", 21856 => "0000000000000000", 21857 => "0000000000000000", 21858 => "0000000000000000", 21859 => "0000000000000000", 21860 => "0000000000000000", 21861 => "0000000000000000", 21862 => "0000000000000000", 21863 => "0000000000000000", 21864 => "0000000000000000", 21865 => "0000000000000000", 21866 => "0000000000000000", 21867 => "0000000000000000", 21868 => "0000000000000000", 21869 => "0000000000000000", 21870 => "0000000000000000", 21871 => "0000000000000000", 21872 => "0000000000000000", 21873 => "0000000000000000", 21874 => "0000000000000000", 21875 => "0000000000000000", 21876 => "0000000000000000", 21877 => "0000000000000000", 21878 => "0000000000000000", 21879 => "0000000000000000", 21880 => "0000000000000000", 21881 => "0000000000000000", 21882 => "0000000000000000", 21883 => "0000000000000000", 21884 => "0000000000000000", 21885 => "0000000000000000", 21886 => "0000000000000000", 21887 => "0000000000000000", 21888 => "0000000000000000", 21889 => "0000000000000000", 21890 => "0000000000000000", 21891 => "0000000000000000", 21892 => "0000000000000000", 21893 => "0000000000000000", 21894 => "0000000000000000", 21895 => "0000000000000000", 21896 => "0000000000000000", 21897 => "0000000000000000", 21898 => "0000000000000000", 21899 => "0000000000000000", 21900 => "0000000000000000", 21901 => "0000000000000000", 21902 => "0000000000000000", 21903 => "0000000000000000", 21904 => "0000000000000000", 21905 => "0000000000000000", 21906 => "0000000000000000", 21907 => "0000000000000000", 21908 => "0000000000000000", 21909 => "0000000000000000", 21910 => "0000000000000000", 21911 => "0000000000000000", 21912 => "0000000000000000", 21913 => "0000000000000000", 21914 => "0000000000000000", 21915 => "0000000000000000", 21916 => "0000000000000000", 21917 => "0000000000000000", 21918 => "0000000000000000", 21919 => "0000000000000000", 21920 => "0000000000000000", 21921 => "0000000000000000", 21922 => "0000000000000000", 21923 => "0000000000000000", 21924 => "0000000000000000", 21925 => "0000000000000000", 21926 => "0000000000000000", 21927 => "0000000000000000", 21928 => "0000000000000000", 21929 => "0000000000000000", 21930 => "0000000000000000", 21931 => "0000000000000000", 21932 => "0000000000000000", 21933 => "0000000000000000", 21934 => "0000000000000000", 21935 => "0000000000000000", 21936 => "0000000000000000", 21937 => "0000000000000000", 21938 => "0000000000000000", 21939 => "0000000000000000", 21940 => "0000000000000000", 21941 => "0000000000000000", 21942 => "0000000000000000", 21943 => "0000000000000000", 21944 => "0000000000000000", 21945 => "0000000000000000", 21946 => "0000000000000000", 21947 => "0000000000000000", 21948 => "0000000000000000", 21949 => "0000000000000000", 21950 => "0000000000000000", 21951 => "0000000000000000", 21952 => "0000000000000000", 21953 => "0000000000000000", 21954 => "0000000000000000", 21955 => "0000000000000000", 21956 => "0000000000000000", 21957 => "0000000000000000", 21958 => "0000000000000000", 21959 => "0000000000000000", 21960 => "0000000000000000", 21961 => "0000000000000000", 21962 => "0000000000000000", 21963 => "0000000000000000", 21964 => "0000000000000000", 21965 => "0000000000000000", 21966 => "0000000000000000", 21967 => "0000000000000000", 21968 => "0000000000000000", 21969 => "0000000000000000", 21970 => "0000000000000000", 21971 => "0000000000000000", 21972 => "0000000000000000", 21973 => "0000000000000000", 21974 => "0000000000000000", 21975 => "0000000000000000", 21976 => "0000000000000000", 21977 => "0000000000000000", 21978 => "0000000000000000", 21979 => "0000000000000000", 21980 => "0000000000000000", 21981 => "0000000000000000", 21982 => "0000000000000000", 21983 => "0000000000000000", 21984 => "0000000000000000", 21985 => "0000000000000000", 21986 => "0000000000000000", 21987 => "0000000000000000", 21988 => "0000000000000000", 21989 => "0000000000000000", 21990 => "0000000000000000", 21991 => "0000000000000000", 21992 => "0000000000000000", 21993 => "0000000000000000", 21994 => "0000000000000000", 21995 => "0000000000000000", 21996 => "0000000000000000", 21997 => "0000000000000000", 21998 => "0000000000000000", 21999 => "0000000000000000", 22000 => "0000000000000000", 22001 => "0000000000000000", 22002 => "0000000000000000", 22003 => "0000000000000000", 22004 => "0000000000000000", 22005 => "0000000000000000", 22006 => "0000000000000000", 22007 => "0000000000000000", 22008 => "0000000000000000", 22009 => "0000000000000000", 22010 => "0000000000000000", 22011 => "0000000000000000", 22012 => "0000000000000000", 22013 => "0000000000000000", 22014 => "0000000000000000", 22015 => "0000000000000000", 22016 => "0000000000000000", 22017 => "0000000000000000", 22018 => "0000000000000000", 22019 => "0000000000000000", 22020 => "0000000000000000", 22021 => "0000000000000000", 22022 => "0000000000000000", 22023 => "0000000000000000", 22024 => "0000000000000000", 22025 => "0000000000000000", 22026 => "0000000000000000", 22027 => "0000000000000000", 22028 => "0000000000000000", 22029 => "0000000000000000", 22030 => "0000000000000000", 22031 => "0000000000000000", 22032 => "0000000000000000", 22033 => "0000000000000000", 22034 => "0000000000000000", 22035 => "0000000000000000", 22036 => "0000000000000000", 22037 => "0000000000000000", 22038 => "0000000000000000", 22039 => "0000000000000000", 22040 => "0000000000000000", 22041 => "0000000000000000", 22042 => "0000000000000000", 22043 => "0000000000000000", 22044 => "0000000000000000", 22045 => "0000000000000000", 22046 => "0000000000000000", 22047 => "0000000000000000", 22048 => "0000000000000000", 22049 => "0000000000000000", 22050 => "0000000000000000", 22051 => "0000000000000000", 22052 => "0000000000000000", 22053 => "0000000000000000", 22054 => "0000000000000000", 22055 => "0000000000000000", 22056 => "0000000000000000", 22057 => "0000000000000000", 22058 => "0000000000000000", 22059 => "0000000000000000", 22060 => "0000000000000000", 22061 => "0000000000000000", 22062 => "0000000000000000", 22063 => "0000000000000000", 22064 => "0000000000000000", 22065 => "0000000000000000", 22066 => "0000000000000000", 22067 => "0000000000000000", 22068 => "0000000000000000", 22069 => "0000000000000000", 22070 => "0000000000000000", 22071 => "0000000000000000", 22072 => "0000000000000000", 22073 => "0000000000000000", 22074 => "0000000000000000", 22075 => "0000000000000000", 22076 => "0000000000000000", 22077 => "0000000000000000", 22078 => "0000000000000000", 22079 => "0000000000000000", 22080 => "0000000000000000", 22081 => "0000000000000000", 22082 => "0000000000000000", 22083 => "0000000000000000", 22084 => "0000000000000000", 22085 => "0000000000000000", 22086 => "0000000000000000", 22087 => "0000000000000000", 22088 => "0000000000000000", 22089 => "0000000000000000", 22090 => "0000000000000000", 22091 => "0000000000000000", 22092 => "0000000000000000", 22093 => "0000000000000000", 22094 => "0000000000000000", 22095 => "0000000000000000", 22096 => "0000000000000000", 22097 => "0000000000000000", 22098 => "0000000000000000", 22099 => "0000000000000000", 22100 => "0000000000000000", 22101 => "0000000000000000", 22102 => "0000000000000000", 22103 => "0000000000000000", 22104 => "0000000000000000", 22105 => "0000000000000000", 22106 => "0000000000000000", 22107 => "0000000000000000", 22108 => "0000000000000000", 22109 => "0000000000000000", 22110 => "0000000000000000", 22111 => "0000000000000000", 22112 => "0000000000000000", 22113 => "0000000000000000", 22114 => "0000000000000000", 22115 => "0000000000000000", 22116 => "0000000000000000", 22117 => "0000000000000000", 22118 => "0000000000000000", 22119 => "0000000000000000", 22120 => "0000000000000000", 22121 => "0000000000000000", 22122 => "0000000000000000", 22123 => "0000000000000000", 22124 => "0000000000000000", 22125 => "0000000000000000", 22126 => "0000000000000000", 22127 => "0000000000000000", 22128 => "0000000000000000", 22129 => "0000000000000000", 22130 => "0000000000000000", 22131 => "0000000000000000", 22132 => "0000000000000000", 22133 => "0000000000000000", 22134 => "0000000000000000", 22135 => "0000000000000000", 22136 => "0000000000000000", 22137 => "0000000000000000", 22138 => "0000000000000000", 22139 => "0000000000000000", 22140 => "0000000000000000", 22141 => "0000000000000000", 22142 => "0000000000000000", 22143 => "0000000000000000", 22144 => "0000000000000000", 22145 => "0000000000000000", 22146 => "0000000000000000", 22147 => "0000000000000000", 22148 => "0000000000000000", 22149 => "0000000000000000", 22150 => "0000000000000000", 22151 => "0000000000000000", 22152 => "0000000000000000", 22153 => "0000000000000000", 22154 => "0000000000000000", 22155 => "0000000000000000", 22156 => "0000000000000000", 22157 => "0000000000000000", 22158 => "0000000000000000", 22159 => "0000000000000000", 22160 => "0000000000000000", 22161 => "0000000000000000", 22162 => "0000000000000000", 22163 => "0000000000000000", 22164 => "0000000000000000", 22165 => "0000000000000000", 22166 => "0000000000000000", 22167 => "0000000000000000", 22168 => "0000000000000000", 22169 => "0000000000000000", 22170 => "0000000000000000", 22171 => "0000000000000000", 22172 => "0000000000000000", 22173 => "0000000000000000", 22174 => "0000000000000000", 22175 => "0000000000000000", 22176 => "0000000000000000", 22177 => "0000000000000000", 22178 => "0000000000000000", 22179 => "0000000000000000", 22180 => "0000000000000000", 22181 => "0000000000000000", 22182 => "0000000000000000", 22183 => "0000000000000000", 22184 => "0000000000000000", 22185 => "0000000000000000", 22186 => "0000000000000000", 22187 => "0000000000000000", 22188 => "0000000000000000", 22189 => "0000000000000000", 22190 => "0000000000000000", 22191 => "0000000000000000", 22192 => "0000000000000000", 22193 => "0000000000000000", 22194 => "0000000000000000", 22195 => "0000000000000000", 22196 => "0000000000000000", 22197 => "0000000000000000", 22198 => "0000000000000000", 22199 => "0000000000000000", 22200 => "0000000000000000", 22201 => "0000000000000000", 22202 => "0000000000000000", 22203 => "0000000000000000", 22204 => "0000000000000000", 22205 => "0000000000000000", 22206 => "0000000000000000", 22207 => "0000000000000000", 22208 => "0000000000000000", 22209 => "0000000000000000", 22210 => "0000000000000000", 22211 => "0000000000000000", 22212 => "0000000000000000", 22213 => "0000000000000000", 22214 => "0000000000000000", 22215 => "0000000000000000", 22216 => "0000000000000000", 22217 => "0000000000000000", 22218 => "0000000000000000", 22219 => "0000000000000000", 22220 => "0000000000000000", 22221 => "0000000000000000", 22222 => "0000000000000000", 22223 => "0000000000000000", 22224 => "0000000000000000", 22225 => "0000000000000000", 22226 => "0000000000000000", 22227 => "0000000000000000", 22228 => "0000000000000000", 22229 => "0000000000000000", 22230 => "0000000000000000", 22231 => "0000000000000000", 22232 => "0000000000000000", 22233 => "0000000000000000", 22234 => "0000000000000000", 22235 => "0000000000000000", 22236 => "0000000000000000", 22237 => "0000000000000000", 22238 => "0000000000000000", 22239 => "0000000000000000", 22240 => "0000000000000000", 22241 => "0000000000000000", 22242 => "0000000000000000", 22243 => "0000000000000000", 22244 => "0000000000000000", 22245 => "0000000000000000", 22246 => "0000000000000000", 22247 => "0000000000000000", 22248 => "0000000000000000", 22249 => "0000000000000000", 22250 => "0000000000000000", 22251 => "0000000000000000", 22252 => "0000000000000000", 22253 => "0000000000000000", 22254 => "0000000000000000", 22255 => "0000000000000000", 22256 => "0000000000000000", 22257 => "0000000000000000", 22258 => "0000000000000000", 22259 => "0000000000000000", 22260 => "0000000000000000", 22261 => "0000000000000000", 22262 => "0000000000000000", 22263 => "0000000000000000", 22264 => "0000000000000000", 22265 => "0000000000000000", 22266 => "0000000000000000", 22267 => "0000000000000000", 22268 => "0000000000000000", 22269 => "0000000000000000", 22270 => "0000000000000000", 22271 => "0000000000000000", 22272 => "0000000000000000", 22273 => "0000000000000000", 22274 => "0000000000000000", 22275 => "0000000000000000", 22276 => "0000000000000000", 22277 => "0000000000000000", 22278 => "0000000000000000", 22279 => "0000000000000000", 22280 => "0000000000000000", 22281 => "0000000000000000", 22282 => "0000000000000000", 22283 => "0000000000000000", 22284 => "0000000000000000", 22285 => "0000000000000000", 22286 => "0000000000000000", 22287 => "0000000000000000", 22288 => "0000000000000000", 22289 => "0000000000000000", 22290 => "0000000000000000", 22291 => "0000000000000000", 22292 => "0000000000000000", 22293 => "0000000000000000", 22294 => "0000000000000000", 22295 => "0000000000000000", 22296 => "0000000000000000", 22297 => "0000000000000000", 22298 => "0000000000000000", 22299 => "0000000000000000", 22300 => "0000000000000000", 22301 => "0000000000000000", 22302 => "0000000000000000", 22303 => "0000000000000000", 22304 => "0000000000000000", 22305 => "0000000000000000", 22306 => "0000000000000000", 22307 => "0000000000000000", 22308 => "0000000000000000", 22309 => "0000000000000000", 22310 => "0000000000000000", 22311 => "0000000000000000", 22312 => "0000000000000000", 22313 => "0000000000000000", 22314 => "0000000000000000", 22315 => "0000000000000000", 22316 => "0000000000000000", 22317 => "0000000000000000", 22318 => "0000000000000000", 22319 => "0000000000000000", 22320 => "0000000000000000", 22321 => "0000000000000000", 22322 => "0000000000000000", 22323 => "0000000000000000", 22324 => "0000000000000000", 22325 => "0000000000000000", 22326 => "0000000000000000", 22327 => "0000000000000000", 22328 => "0000000000000000", 22329 => "0000000000000000", 22330 => "0000000000000000", 22331 => "0000000000000000", 22332 => "0000000000000000", 22333 => "0000000000000000", 22334 => "0000000000000000", 22335 => "0000000000000000", 22336 => "0000000000000000", 22337 => "0000000000000000", 22338 => "0000000000000000", 22339 => "0000000000000000", 22340 => "0000000000000000", 22341 => "0000000000000000", 22342 => "0000000000000000", 22343 => "0000000000000000", 22344 => "0000000000000000", 22345 => "0000000000000000", 22346 => "0000000000000000", 22347 => "0000000000000000", 22348 => "0000000000000000", 22349 => "0000000000000000", 22350 => "0000000000000000", 22351 => "0000000000000000", 22352 => "0000000000000000", 22353 => "0000000000000000", 22354 => "0000000000000000", 22355 => "0000000000000000", 22356 => "0000000000000000", 22357 => "0000000000000000", 22358 => "0000000000000000", 22359 => "0000000000000000", 22360 => "0000000000000000", 22361 => "0000000000000000", 22362 => "0000000000000000", 22363 => "0000000000000000", 22364 => "0000000000000000", 22365 => "0000000000000000", 22366 => "0000000000000000", 22367 => "0000000000000000", 22368 => "0000000000000000", 22369 => "0000000000000000", 22370 => "0000000000000000", 22371 => "0000000000000000", 22372 => "0000000000000000", 22373 => "0000000000000000", 22374 => "0000000000000000", 22375 => "0000000000000000", 22376 => "0000000000000000", 22377 => "0000000000000000", 22378 => "0000000000000000", 22379 => "0000000000000000", 22380 => "0000000000000000", 22381 => "0000000000000000", 22382 => "0000000000000000", 22383 => "0000000000000000", 22384 => "0000000000000000", 22385 => "0000000000000000", 22386 => "0000000000000000", 22387 => "0000000000000000", 22388 => "0000000000000000", 22389 => "0000000000000000", 22390 => "0000000000000000", 22391 => "0000000000000000", 22392 => "0000000000000000", 22393 => "0000000000000000", 22394 => "0000000000000000", 22395 => "0000000000000000", 22396 => "0000000000000000", 22397 => "0000000000000000", 22398 => "0000000000000000", 22399 => "0000000000000000", 22400 => "0000000000000000", 22401 => "0000000000000000", 22402 => "0000000000000000", 22403 => "0000000000000000", 22404 => "0000000000000000", 22405 => "0000000000000000", 22406 => "0000000000000000", 22407 => "0000000000000000", 22408 => "0000000000000000", 22409 => "0000000000000000", 22410 => "0000000000000000", 22411 => "0000000000000000", 22412 => "0000000000000000", 22413 => "0000000000000000", 22414 => "0000000000000000", 22415 => "0000000000000000", 22416 => "0000000000000000", 22417 => "0000000000000000", 22418 => "0000000000000000", 22419 => "0000000000000000", 22420 => "0000000000000000", 22421 => "0000000000000000", 22422 => "0000000000000000", 22423 => "0000000000000000", 22424 => "0000000000000000", 22425 => "0000000000000000", 22426 => "0000000000000000", 22427 => "0000000000000000", 22428 => "0000000000000000", 22429 => "0000000000000000", 22430 => "0000000000000000", 22431 => "0000000000000000", 22432 => "0000000000000000", 22433 => "0000000000000000", 22434 => "0000000000000000", 22435 => "0000000000000000", 22436 => "0000000000000000", 22437 => "0000000000000000", 22438 => "0000000000000000", 22439 => "0000000000000000", 22440 => "0000000000000000", 22441 => "0000000000000000", 22442 => "0000000000000000", 22443 => "0000000000000000", 22444 => "0000000000000000", 22445 => "0000000000000000", 22446 => "0000000000000000", 22447 => "0000000000000000", 22448 => "0000000000000000", 22449 => "0000000000000000", 22450 => "0000000000000000", 22451 => "0000000000000000", 22452 => "0000000000000000", 22453 => "0000000000000000", 22454 => "0000000000000000", 22455 => "0000000000000000", 22456 => "0000000000000000", 22457 => "0000000000000000", 22458 => "0000000000000000", 22459 => "0000000000000000", 22460 => "0000000000000000", 22461 => "0000000000000000", 22462 => "0000000000000000", 22463 => "0000000000000000", 22464 => "0000000000000000", 22465 => "0000000000000000", 22466 => "0000000000000000", 22467 => "0000000000000000", 22468 => "0000000000000000", 22469 => "0000000000000000", 22470 => "0000000000000000", 22471 => "0000000000000000", 22472 => "0000000000000000", 22473 => "0000000000000000", 22474 => "0000000000000000", 22475 => "0000000000000000", 22476 => "0000000000000000", 22477 => "0000000000000000", 22478 => "0000000000000000", 22479 => "0000000000000000", 22480 => "0000000000000000", 22481 => "0000000000000000", 22482 => "0000000000000000", 22483 => "0000000000000000", 22484 => "0000000000000000", 22485 => "0000000000000000", 22486 => "0000000000000000", 22487 => "0000000000000000", 22488 => "0000000000000000", 22489 => "0000000000000000", 22490 => "0000000000000000", 22491 => "0000000000000000", 22492 => "0000000000000000", 22493 => "0000000000000000", 22494 => "0000000000000000", 22495 => "0000000000000000", 22496 => "0000000000000000", 22497 => "0000000000000000", 22498 => "0000000000000000", 22499 => "0000000000000000", 22500 => "0000000000000000", 22501 => "0000000000000000", 22502 => "0000000000000000", 22503 => "0000000000000000", 22504 => "0000000000000000", 22505 => "0000000000000000", 22506 => "0000000000000000", 22507 => "0000000000000000", 22508 => "0000000000000000", 22509 => "0000000000000000", 22510 => "0000000000000000", 22511 => "0000000000000000", 22512 => "0000000000000000", 22513 => "0000000000000000", 22514 => "0000000000000000", 22515 => "0000000000000000", 22516 => "0000000000000000", 22517 => "0000000000000000", 22518 => "0000000000000000", 22519 => "0000000000000000", 22520 => "0000000000000000", 22521 => "0000000000000000", 22522 => "0000000000000000", 22523 => "0000000000000000", 22524 => "0000000000000000", 22525 => "0000000000000000", 22526 => "0000000000000000", 22527 => "0000000000000000", 22528 => "0000000000000000", 22529 => "0000000000000000", 22530 => "0000000000000000", 22531 => "0000000000000000", 22532 => "0000000000000000", 22533 => "0000000000000000", 22534 => "0000000000000000", 22535 => "0000000000000000", 22536 => "0000000000000000", 22537 => "0000000000000000", 22538 => "0000000000000000", 22539 => "0000000000000000", 22540 => "0000000000000000", 22541 => "0000000000000000", 22542 => "0000000000000000", 22543 => "0000000000000000", 22544 => "0000000000000000", 22545 => "0000000000000000", 22546 => "0000000000000000", 22547 => "0000000000000000", 22548 => "0000000000000000", 22549 => "0000000000000000", 22550 => "0000000000000000", 22551 => "0000000000000000", 22552 => "0000000000000000", 22553 => "0000000000000000", 22554 => "0000000000000000", 22555 => "0000000000000000", 22556 => "0000000000000000", 22557 => "0000000000000000", 22558 => "0000000000000000", 22559 => "0000000000000000", 22560 => "0000000000000000", 22561 => "0000000000000000", 22562 => "0000000000000000", 22563 => "0000000000000000", 22564 => "0000000000000000", 22565 => "0000000000000000", 22566 => "0000000000000000", 22567 => "0000000000000000", 22568 => "0000000000000000", 22569 => "0000000000000000", 22570 => "0000000000000000", 22571 => "0000000000000000", 22572 => "0000000000000000", 22573 => "0000000000000000", 22574 => "0000000000000000", 22575 => "0000000000000000", 22576 => "0000000000000000", 22577 => "0000000000000000", 22578 => "0000000000000000", 22579 => "0000000000000000", 22580 => "0000000000000000", 22581 => "0000000000000000", 22582 => "0000000000000000", 22583 => "0000000000000000", 22584 => "0000000000000000", 22585 => "0000000000000000", 22586 => "0000000000000000", 22587 => "0000000000000000", 22588 => "0000000000000000", 22589 => "0000000000000000", 22590 => "0000000000000000", 22591 => "0000000000000000", 22592 => "0000000000000000", 22593 => "0000000000000000", 22594 => "0000000000000000", 22595 => "0000000000000000", 22596 => "0000000000000000", 22597 => "0000000000000000", 22598 => "0000000000000000", 22599 => "0000000000000000", 22600 => "0000000000000000", 22601 => "0000000000000000", 22602 => "0000000000000000", 22603 => "0000000000000000", 22604 => "0000000000000000", 22605 => "0000000000000000", 22606 => "0000000000000000", 22607 => "0000000000000000", 22608 => "0000000000000000", 22609 => "0000000000000000", 22610 => "0000000000000000", 22611 => "0000000000000000", 22612 => "0000000000000000", 22613 => "0000000000000000", 22614 => "0000000000000000", 22615 => "0000000000000000", 22616 => "0000000000000000", 22617 => "0000000000000000", 22618 => "0000000000000000", 22619 => "0000000000000000", 22620 => "0000000000000000", 22621 => "0000000000000000", 22622 => "0000000000000000", 22623 => "0000000000000000", 22624 => "0000000000000000", 22625 => "0000000000000000", 22626 => "0000000000000000", 22627 => "0000000000000000", 22628 => "0000000000000000", 22629 => "0000000000000000", 22630 => "0000000000000000", 22631 => "0000000000000000", 22632 => "0000000000000000", 22633 => "0000000000000000", 22634 => "0000000000000000", 22635 => "0000000000000000", 22636 => "0000000000000000", 22637 => "0000000000000000", 22638 => "0000000000000000", 22639 => "0000000000000000", 22640 => "0000000000000000", 22641 => "0000000000000000", 22642 => "0000000000000000", 22643 => "0000000000000000", 22644 => "0000000000000000", 22645 => "0000000000000000", 22646 => "0000000000000000", 22647 => "0000000000000000", 22648 => "0000000000000000", 22649 => "0000000000000000", 22650 => "0000000000000000", 22651 => "0000000000000000", 22652 => "0000000000000000", 22653 => "0000000000000000", 22654 => "0000000000000000", 22655 => "0000000000000000", 22656 => "0000000000000000", 22657 => "0000000000000000", 22658 => "0000000000000000", 22659 => "0000000000000000", 22660 => "0000000000000000", 22661 => "0000000000000000", 22662 => "0000000000000000", 22663 => "0000000000000000", 22664 => "0000000000000000", 22665 => "0000000000000000", 22666 => "0000000000000000", 22667 => "0000000000000000", 22668 => "0000000000000000", 22669 => "0000000000000000", 22670 => "0000000000000000", 22671 => "0000000000000000", 22672 => "0000000000000000", 22673 => "0000000000000000", 22674 => "0000000000000000", 22675 => "0000000000000000", 22676 => "0000000000000000", 22677 => "0000000000000000", 22678 => "0000000000000000", 22679 => "0000000000000000", 22680 => "0000000000000000", 22681 => "0000000000000000", 22682 => "0000000000000000", 22683 => "0000000000000000", 22684 => "0000000000000000", 22685 => "0000000000000000", 22686 => "0000000000000000", 22687 => "0000000000000000", 22688 => "0000000000000000", 22689 => "0000000000000000", 22690 => "0000000000000000", 22691 => "0000000000000000", 22692 => "0000000000000000", 22693 => "0000000000000000", 22694 => "0000000000000000", 22695 => "0000000000000000", 22696 => "0000000000000000", 22697 => "0000000000000000", 22698 => "0000000000000000", 22699 => "0000000000000000", 22700 => "0000000000000000", 22701 => "0000000000000000", 22702 => "0000000000000000", 22703 => "0000000000000000", 22704 => "0000000000000000", 22705 => "0000000000000000", 22706 => "0000000000000000", 22707 => "0000000000000000", 22708 => "0000000000000000", 22709 => "0000000000000000", 22710 => "0000000000000000", 22711 => "0000000000000000", 22712 => "0000000000000000", 22713 => "0000000000000000", 22714 => "0000000000000000", 22715 => "0000000000000000", 22716 => "0000000000000000", 22717 => "0000000000000000", 22718 => "0000000000000000", 22719 => "0000000000000000", 22720 => "0000000000000000", 22721 => "0000000000000000", 22722 => "0000000000000000", 22723 => "0000000000000000", 22724 => "0000000000000000", 22725 => "0000000000000000", 22726 => "0000000000000000", 22727 => "0000000000000000", 22728 => "0000000000000000", 22729 => "0000000000000000", 22730 => "0000000000000000", 22731 => "0000000000000000", 22732 => "0000000000000000", 22733 => "0000000000000000", 22734 => "0000000000000000", 22735 => "0000000000000000", 22736 => "0000000000000000", 22737 => "0000000000000000", 22738 => "0000000000000000", 22739 => "0000000000000000", 22740 => "0000000000000000", 22741 => "0000000000000000", 22742 => "0000000000000000", 22743 => "0000000000000000", 22744 => "0000000000000000", 22745 => "0000000000000000", 22746 => "0000000000000000", 22747 => "0000000000000000", 22748 => "0000000000000000", 22749 => "0000000000000000", 22750 => "0000000000000000", 22751 => "0000000000000000", 22752 => "0000000000000000", 22753 => "0000000000000000", 22754 => "0000000000000000", 22755 => "0000000000000000", 22756 => "0000000000000000", 22757 => "0000000000000000", 22758 => "0000000000000000", 22759 => "0000000000000000", 22760 => "0000000000000000", 22761 => "0000000000000000", 22762 => "0000000000000000", 22763 => "0000000000000000", 22764 => "0000000000000000", 22765 => "0000000000000000", 22766 => "0000000000000000", 22767 => "0000000000000000", 22768 => "0000000000000000", 22769 => "0000000000000000", 22770 => "0000000000000000", 22771 => "0000000000000000", 22772 => "0000000000000000", 22773 => "0000000000000000", 22774 => "0000000000000000", 22775 => "0000000000000000", 22776 => "0000000000000000", 22777 => "0000000000000000", 22778 => "0000000000000000", 22779 => "0000000000000000", 22780 => "0000000000000000", 22781 => "0000000000000000", 22782 => "0000000000000000", 22783 => "0000000000000000", 22784 => "0000000000000000", 22785 => "0000000000000000", 22786 => "0000000000000000", 22787 => "0000000000000000", 22788 => "0000000000000000", 22789 => "0000000000000000", 22790 => "0000000000000000", 22791 => "0000000000000000", 22792 => "0000000000000000", 22793 => "0000000000000000", 22794 => "0000000000000000", 22795 => "0000000000000000", 22796 => "0000000000000000", 22797 => "0000000000000000", 22798 => "0000000000000000", 22799 => "0000000000000000", 22800 => "0000000000000000", 22801 => "0000000000000000", 22802 => "0000000000000000", 22803 => "0000000000000000", 22804 => "0000000000000000", 22805 => "0000000000000000", 22806 => "0000000000000000", 22807 => "0000000000000000", 22808 => "0000000000000000", 22809 => "0000000000000000", 22810 => "0000000000000000", 22811 => "0000000000000000", 22812 => "0000000000000000", 22813 => "0000000000000000", 22814 => "0000000000000000", 22815 => "0000000000000000", 22816 => "0000000000000000", 22817 => "0000000000000000", 22818 => "0000000000000000", 22819 => "0000000000000000", 22820 => "0000000000000000", 22821 => "0000000000000000", 22822 => "0000000000000000", 22823 => "0000000000000000", 22824 => "0000000000000000", 22825 => "0000000000000000", 22826 => "0000000000000000", 22827 => "0000000000000000", 22828 => "0000000000000000", 22829 => "0000000000000000", 22830 => "0000000000000000", 22831 => "0000000000000000", 22832 => "0000000000000000", 22833 => "0000000000000000", 22834 => "0000000000000000", 22835 => "0000000000000000", 22836 => "0000000000000000", 22837 => "0000000000000000", 22838 => "0000000000000000", 22839 => "0000000000000000", 22840 => "0000000000000000", 22841 => "0000000000000000", 22842 => "0000000000000000", 22843 => "0000000000000000", 22844 => "0000000000000000", 22845 => "0000000000000000", 22846 => "0000000000000000", 22847 => "0000000000000000", 22848 => "0000000000000000", 22849 => "0000000000000000", 22850 => "0000000000000000", 22851 => "0000000000000000", 22852 => "0000000000000000", 22853 => "0000000000000000", 22854 => "0000000000000000", 22855 => "0000000000000000", 22856 => "0000000000000000", 22857 => "0000000000000000", 22858 => "0000000000000000", 22859 => "0000000000000000", 22860 => "0000000000000000", 22861 => "0000000000000000", 22862 => "0000000000000000", 22863 => "0000000000000000", 22864 => "0000000000000000", 22865 => "0000000000000000", 22866 => "0000000000000000", 22867 => "0000000000000000", 22868 => "0000000000000000", 22869 => "0000000000000000", 22870 => "0000000000000000", 22871 => "0000000000000000", 22872 => "0000000000000000", 22873 => "0000000000000000", 22874 => "0000000000000000", 22875 => "0000000000000000", 22876 => "0000000000000000", 22877 => "0000000000000000", 22878 => "0000000000000000", 22879 => "0000000000000000", 22880 => "0000000000000000", 22881 => "0000000000000000", 22882 => "0000000000000000", 22883 => "0000000000000000", 22884 => "0000000000000000", 22885 => "0000000000000000", 22886 => "0000000000000000", 22887 => "0000000000000000", 22888 => "0000000000000000", 22889 => "0000000000000000", 22890 => "0000000000000000", 22891 => "0000000000000000", 22892 => "0000000000000000", 22893 => "0000000000000000", 22894 => "0000000000000000", 22895 => "0000000000000000", 22896 => "0000000000000000", 22897 => "0000000000000000", 22898 => "0000000000000000", 22899 => "0000000000000000", 22900 => "0000000000000000", 22901 => "0000000000000000", 22902 => "0000000000000000", 22903 => "0000000000000000", 22904 => "0000000000000000", 22905 => "0000000000000000", 22906 => "0000000000000000", 22907 => "0000000000000000", 22908 => "0000000000000000", 22909 => "0000000000000000", 22910 => "0000000000000000", 22911 => "0000000000000000", 22912 => "0000000000000000", 22913 => "0000000000000000", 22914 => "0000000000000000", 22915 => "0000000000000000", 22916 => "0000000000000000", 22917 => "0000000000000000", 22918 => "0000000000000000", 22919 => "0000000000000000", 22920 => "0000000000000000", 22921 => "0000000000000000", 22922 => "0000000000000000", 22923 => "0000000000000000", 22924 => "0000000000000000", 22925 => "0000000000000000", 22926 => "0000000000000000", 22927 => "0000000000000000", 22928 => "0000000000000000", 22929 => "0000000000000000", 22930 => "0000000000000000", 22931 => "0000000000000000", 22932 => "0000000000000000", 22933 => "0000000000000000", 22934 => "0000000000000000", 22935 => "0000000000000000", 22936 => "0000000000000000", 22937 => "0000000000000000", 22938 => "0000000000000000", 22939 => "0000000000000000", 22940 => "0000000000000000", 22941 => "0000000000000000", 22942 => "0000000000000000", 22943 => "0000000000000000", 22944 => "0000000000000000", 22945 => "0000000000000000", 22946 => "0000000000000000", 22947 => "0000000000000000", 22948 => "0000000000000000", 22949 => "0000000000000000", 22950 => "0000000000000000", 22951 => "0000000000000000", 22952 => "0000000000000000", 22953 => "0000000000000000", 22954 => "0000000000000000", 22955 => "0000000000000000", 22956 => "0000000000000000", 22957 => "0000000000000000", 22958 => "0000000000000000", 22959 => "0000000000000000", 22960 => "0000000000000000", 22961 => "0000000000000000", 22962 => "0000000000000000", 22963 => "0000000000000000", 22964 => "0000000000000000", 22965 => "0000000000000000", 22966 => "0000000000000000", 22967 => "0000000000000000", 22968 => "0000000000000000", 22969 => "0000000000000000", 22970 => "0000000000000000", 22971 => "0000000000000000", 22972 => "0000000000000000", 22973 => "0000000000000000", 22974 => "0000000000000000", 22975 => "0000000000000000", 22976 => "0000000000000000", 22977 => "0000000000000000", 22978 => "0000000000000000", 22979 => "0000000000000000", 22980 => "0000000000000000", 22981 => "0000000000000000", 22982 => "0000000000000000", 22983 => "0000000000000000", 22984 => "0000000000000000", 22985 => "0000000000000000", 22986 => "0000000000000000", 22987 => "0000000000000000", 22988 => "0000000000000000", 22989 => "0000000000000000", 22990 => "0000000000000000", 22991 => "0000000000000000", 22992 => "0000000000000000", 22993 => "0000000000000000", 22994 => "0000000000000000", 22995 => "0000000000000000", 22996 => "0000000000000000", 22997 => "0000000000000000", 22998 => "0000000000000000", 22999 => "0000000000000000", 23000 => "0000000000000000", 23001 => "0000000000000000", 23002 => "0000000000000000", 23003 => "0000000000000000", 23004 => "0000000000000000", 23005 => "0000000000000000", 23006 => "0000000000000000", 23007 => "0000000000000000", 23008 => "0000000000000000", 23009 => "0000000000000000", 23010 => "0000000000000000", 23011 => "0000000000000000", 23012 => "0000000000000000", 23013 => "0000000000000000", 23014 => "0000000000000000", 23015 => "0000000000000000", 23016 => "0000000000000000", 23017 => "0000000000000000", 23018 => "0000000000000000", 23019 => "0000000000000000", 23020 => "0000000000000000", 23021 => "0000000000000000", 23022 => "0000000000000000", 23023 => "0000000000000000", 23024 => "0000000000000000", 23025 => "0000000000000000", 23026 => "0000000000000000", 23027 => "0000000000000000", 23028 => "0000000000000000", 23029 => "0000000000000000", 23030 => "0000000000000000", 23031 => "0000000000000000", 23032 => "0000000000000000", 23033 => "0000000000000000", 23034 => "0000000000000000", 23035 => "0000000000000000", 23036 => "0000000000000000", 23037 => "0000000000000000", 23038 => "0000000000000000", 23039 => "0000000000000000", 23040 => "0000000000000000", 23041 => "0000000000000000", 23042 => "0000000000000000", 23043 => "0000000000000000", 23044 => "0000000000000000", 23045 => "0000000000000000", 23046 => "0000000000000000", 23047 => "0000000000000000", 23048 => "0000000000000000", 23049 => "0000000000000000", 23050 => "0000000000000000", 23051 => "0000000000000000", 23052 => "0000000000000000", 23053 => "0000000000000000", 23054 => "0000000000000000", 23055 => "0000000000000000", 23056 => "0000000000000000", 23057 => "0000000000000000", 23058 => "0000000000000000", 23059 => "0000000000000000", 23060 => "0000000000000000", 23061 => "0000000000000000", 23062 => "0000000000000000", 23063 => "0000000000000000", 23064 => "0000000000000000", 23065 => "0000000000000000", 23066 => "0000000000000000", 23067 => "0000000000000000", 23068 => "0000000000000000", 23069 => "0000000000000000", 23070 => "0000000000000000", 23071 => "0000000000000000", 23072 => "0000000000000000", 23073 => "0000000000000000", 23074 => "0000000000000000", 23075 => "0000000000000000", 23076 => "0000000000000000", 23077 => "0000000000000000", 23078 => "0000000000000000", 23079 => "0000000000000000", 23080 => "0000000000000000", 23081 => "0000000000000000", 23082 => "0000000000000000", 23083 => "0000000000000000", 23084 => "0000000000000000", 23085 => "0000000000000000", 23086 => "0000000000000000", 23087 => "0000000000000000", 23088 => "0000000000000000", 23089 => "0000000000000000", 23090 => "0000000000000000", 23091 => "0000000000000000", 23092 => "0000000000000000", 23093 => "0000000000000000", 23094 => "0000000000000000", 23095 => "0000000000000000", 23096 => "0000000000000000", 23097 => "0000000000000000", 23098 => "0000000000000000", 23099 => "0000000000000000", 23100 => "0000000000000000", 23101 => "0000000000000000", 23102 => "0000000000000000", 23103 => "0000000000000000", 23104 => "0000000000000000", 23105 => "0000000000000000", 23106 => "0000000000000000", 23107 => "0000000000000000", 23108 => "0000000000000000", 23109 => "0000000000000000", 23110 => "0000000000000000", 23111 => "0000000000000000", 23112 => "0000000000000000", 23113 => "0000000000000000", 23114 => "0000000000000000", 23115 => "0000000000000000", 23116 => "0000000000000000", 23117 => "0000000000000000", 23118 => "0000000000000000", 23119 => "0000000000000000", 23120 => "0000000000000000", 23121 => "0000000000000000", 23122 => "0000000000000000", 23123 => "0000000000000000", 23124 => "0000000000000000", 23125 => "0000000000000000", 23126 => "0000000000000000", 23127 => "0000000000000000", 23128 => "0000000000000000", 23129 => "0000000000000000", 23130 => "0000000000000000", 23131 => "0000000000000000", 23132 => "0000000000000000", 23133 => "0000000000000000", 23134 => "0000000000000000", 23135 => "0000000000000000", 23136 => "0000000000000000", 23137 => "0000000000000000", 23138 => "0000000000000000", 23139 => "0000000000000000", 23140 => "0000000000000000", 23141 => "0000000000000000", 23142 => "0000000000000000", 23143 => "0000000000000000", 23144 => "0000000000000000", 23145 => "0000000000000000", 23146 => "0000000000000000", 23147 => "0000000000000000", 23148 => "0000000000000000", 23149 => "0000000000000000", 23150 => "0000000000000000", 23151 => "0000000000000000", 23152 => "0000000000000000", 23153 => "0000000000000000", 23154 => "0000000000000000", 23155 => "0000000000000000", 23156 => "0000000000000000", 23157 => "0000000000000000", 23158 => "0000000000000000", 23159 => "0000000000000000", 23160 => "0000000000000000", 23161 => "0000000000000000", 23162 => "0000000000000000", 23163 => "0000000000000000", 23164 => "0000000000000000", 23165 => "0000000000000000", 23166 => "0000000000000000", 23167 => "0000000000000000", 23168 => "0000000000000000", 23169 => "0000000000000000", 23170 => "0000000000000000", 23171 => "0000000000000000", 23172 => "0000000000000000", 23173 => "0000000000000000", 23174 => "0000000000000000", 23175 => "0000000000000000", 23176 => "0000000000000000", 23177 => "0000000000000000", 23178 => "0000000000000000", 23179 => "0000000000000000", 23180 => "0000000000000000", 23181 => "0000000000000000", 23182 => "0000000000000000", 23183 => "0000000000000000", 23184 => "0000000000000000", 23185 => "0000000000000000", 23186 => "0000000000000000", 23187 => "0000000000000000", 23188 => "0000000000000000", 23189 => "0000000000000000", 23190 => "0000000000000000", 23191 => "0000000000000000", 23192 => "0000000000000000", 23193 => "0000000000000000", 23194 => "0000000000000000", 23195 => "0000000000000000", 23196 => "0000000000000000", 23197 => "0000000000000000", 23198 => "0000000000000000", 23199 => "0000000000000000", 23200 => "0000000000000000", 23201 => "0000000000000000", 23202 => "0000000000000000", 23203 => "0000000000000000", 23204 => "0000000000000000", 23205 => "0000000000000000", 23206 => "0000000000000000", 23207 => "0000000000000000", 23208 => "0000000000000000", 23209 => "0000000000000000", 23210 => "0000000000000000", 23211 => "0000000000000000", 23212 => "0000000000000000", 23213 => "0000000000000000", 23214 => "0000000000000000", 23215 => "0000000000000000", 23216 => "0000000000000000", 23217 => "0000000000000000", 23218 => "0000000000000000", 23219 => "0000000000000000", 23220 => "0000000000000000", 23221 => "0000000000000000", 23222 => "0000000000000000", 23223 => "0000000000000000", 23224 => "0000000000000000", 23225 => "0000000000000000", 23226 => "0000000000000000", 23227 => "0000000000000000", 23228 => "0000000000000000", 23229 => "0000000000000000", 23230 => "0000000000000000", 23231 => "0000000000000000", 23232 => "0000000000000000", 23233 => "0000000000000000", 23234 => "0000000000000000", 23235 => "0000000000000000", 23236 => "0000000000000000", 23237 => "0000000000000000", 23238 => "0000000000000000", 23239 => "0000000000000000", 23240 => "0000000000000000", 23241 => "0000000000000000", 23242 => "0000000000000000", 23243 => "0000000000000000", 23244 => "0000000000000000", 23245 => "0000000000000000", 23246 => "0000000000000000", 23247 => "0000000000000000", 23248 => "0000000000000000", 23249 => "0000000000000000", 23250 => "0000000000000000", 23251 => "0000000000000000", 23252 => "0000000000000000", 23253 => "0000000000000000", 23254 => "0000000000000000", 23255 => "0000000000000000", 23256 => "0000000000000000", 23257 => "0000000000000000", 23258 => "0000000000000000", 23259 => "0000000000000000", 23260 => "0000000000000000", 23261 => "0000000000000000", 23262 => "0000000000000000", 23263 => "0000000000000000", 23264 => "0000000000000000", 23265 => "0000000000000000", 23266 => "0000000000000000", 23267 => "0000000000000000", 23268 => "0000000000000000", 23269 => "0000000000000000", 23270 => "0000000000000000", 23271 => "0000000000000000", 23272 => "0000000000000000", 23273 => "0000000000000000", 23274 => "0000000000000000", 23275 => "0000000000000000", 23276 => "0000000000000000", 23277 => "0000000000000000", 23278 => "0000000000000000", 23279 => "0000000000000000", 23280 => "0000000000000000", 23281 => "0000000000000000", 23282 => "0000000000000000", 23283 => "0000000000000000", 23284 => "0000000000000000", 23285 => "0000000000000000", 23286 => "0000000000000000", 23287 => "0000000000000000", 23288 => "0000000000000000", 23289 => "0000000000000000", 23290 => "0000000000000000", 23291 => "0000000000000000", 23292 => "0000000000000000", 23293 => "0000000000000000", 23294 => "0000000000000000", 23295 => "0000000000000000", 23296 => "0000000000000000", 23297 => "0000000000000000", 23298 => "0000000000000000", 23299 => "0000000000000000", 23300 => "0000000000000000", 23301 => "0000000000000000", 23302 => "0000000000000000", 23303 => "0000000000000000", 23304 => "0000000000000000", 23305 => "0000000000000000", 23306 => "0000000000000000", 23307 => "0000000000000000", 23308 => "0000000000000000", 23309 => "0000000000000000", 23310 => "0000000000000000", 23311 => "0000000000000000", 23312 => "0000000000000000", 23313 => "0000000000000000", 23314 => "0000000000000000", 23315 => "0000000000000000", 23316 => "0000000000000000", 23317 => "0000000000000000", 23318 => "0000000000000000", 23319 => "0000000000000000", 23320 => "0000000000000000", 23321 => "0000000000000000", 23322 => "0000000000000000", 23323 => "0000000000000000", 23324 => "0000000000000000", 23325 => "0000000000000000", 23326 => "0000000000000000", 23327 => "0000000000000000", 23328 => "0000000000000000", 23329 => "0000000000000000", 23330 => "0000000000000000", 23331 => "0000000000000000", 23332 => "0000000000000000", 23333 => "0000000000000000", 23334 => "0000000000000000", 23335 => "0000000000000000", 23336 => "0000000000000000", 23337 => "0000000000000000", 23338 => "0000000000000000", 23339 => "0000000000000000", 23340 => "0000000000000000", 23341 => "0000000000000000", 23342 => "0000000000000000", 23343 => "0000000000000000", 23344 => "0000000000000000", 23345 => "0000000000000000", 23346 => "0000000000000000", 23347 => "0000000000000000", 23348 => "0000000000000000", 23349 => "0000000000000000", 23350 => "0000000000000000", 23351 => "0000000000000000", 23352 => "0000000000000000", 23353 => "0000000000000000", 23354 => "0000000000000000", 23355 => "0000000000000000", 23356 => "0000000000000000", 23357 => "0000000000000000", 23358 => "0000000000000000", 23359 => "0000000000000000", 23360 => "0000000000000000", 23361 => "0000000000000000", 23362 => "0000000000000000", 23363 => "0000000000000000", 23364 => "0000000000000000", 23365 => "0000000000000000", 23366 => "0000000000000000", 23367 => "0000000000000000", 23368 => "0000000000000000", 23369 => "0000000000000000", 23370 => "0000000000000000", 23371 => "0000000000000000", 23372 => "0000000000000000", 23373 => "0000000000000000", 23374 => "0000000000000000", 23375 => "0000000000000000", 23376 => "0000000000000000", 23377 => "0000000000000000", 23378 => "0000000000000000", 23379 => "0000000000000000", 23380 => "0000000000000000", 23381 => "0000000000000000", 23382 => "0000000000000000", 23383 => "0000000000000000", 23384 => "0000000000000000", 23385 => "0000000000000000", 23386 => "0000000000000000", 23387 => "0000000000000000", 23388 => "0000000000000000", 23389 => "0000000000000000", 23390 => "0000000000000000", 23391 => "0000000000000000", 23392 => "0000000000000000", 23393 => "0000000000000000", 23394 => "0000000000000000", 23395 => "0000000000000000", 23396 => "0000000000000000", 23397 => "0000000000000000", 23398 => "0000000000000000", 23399 => "0000000000000000", 23400 => "0000000000000000", 23401 => "0000000000000000", 23402 => "0000000000000000", 23403 => "0000000000000000", 23404 => "0000000000000000", 23405 => "0000000000000000", 23406 => "0000000000000000", 23407 => "0000000000000000", 23408 => "0000000000000000", 23409 => "0000000000000000", 23410 => "0000000000000000", 23411 => "0000000000000000", 23412 => "0000000000000000", 23413 => "0000000000000000", 23414 => "0000000000000000", 23415 => "0000000000000000", 23416 => "0000000000000000", 23417 => "0000000000000000", 23418 => "0000000000000000", 23419 => "0000000000000000", 23420 => "0000000000000000", 23421 => "0000000000000000", 23422 => "0000000000000000", 23423 => "0000000000000000", 23424 => "0000000000000000", 23425 => "0000000000000000", 23426 => "0000000000000000", 23427 => "0000000000000000", 23428 => "0000000000000000", 23429 => "0000000000000000", 23430 => "0000000000000000", 23431 => "0000000000000000", 23432 => "0000000000000000", 23433 => "0000000000000000", 23434 => "0000000000000000", 23435 => "0000000000000000", 23436 => "0000000000000000", 23437 => "0000000000000000", 23438 => "0000000000000000", 23439 => "0000000000000000", 23440 => "0000000000000000", 23441 => "0000000000000000", 23442 => "0000000000000000", 23443 => "0000000000000000", 23444 => "0000000000000000", 23445 => "0000000000000000", 23446 => "0000000000000000", 23447 => "0000000000000000", 23448 => "0000000000000000", 23449 => "0000000000000000", 23450 => "0000000000000000", 23451 => "0000000000000000", 23452 => "0000000000000000", 23453 => "0000000000000000", 23454 => "0000000000000000", 23455 => "0000000000000000", 23456 => "0000000000000000", 23457 => "0000000000000000", 23458 => "0000000000000000", 23459 => "0000000000000000", 23460 => "0000000000000000", 23461 => "0000000000000000", 23462 => "0000000000000000", 23463 => "0000000000000000", 23464 => "0000000000000000", 23465 => "0000000000000000", 23466 => "0000000000000000", 23467 => "0000000000000000", 23468 => "0000000000000000", 23469 => "0000000000000000", 23470 => "0000000000000000", 23471 => "0000000000000000", 23472 => "0000000000000000", 23473 => "0000000000000000", 23474 => "0000000000000000", 23475 => "0000000000000000", 23476 => "0000000000000000", 23477 => "0000000000000000", 23478 => "0000000000000000", 23479 => "0000000000000000", 23480 => "0000000000000000", 23481 => "0000000000000000", 23482 => "0000000000000000", 23483 => "0000000000000000", 23484 => "0000000000000000", 23485 => "0000000000000000", 23486 => "0000000000000000", 23487 => "0000000000000000", 23488 => "0000000000000000", 23489 => "0000000000000000", 23490 => "0000000000000000", 23491 => "0000000000000000", 23492 => "0000000000000000", 23493 => "0000000000000000", 23494 => "0000000000000000", 23495 => "0000000000000000", 23496 => "0000000000000000", 23497 => "0000000000000000", 23498 => "0000000000000000", 23499 => "0000000000000000", 23500 => "0000000000000000", 23501 => "0000000000000000", 23502 => "0000000000000000", 23503 => "0000000000000000", 23504 => "0000000000000000", 23505 => "0000000000000000", 23506 => "0000000000000000", 23507 => "0000000000000000", 23508 => "0000000000000000", 23509 => "0000000000000000", 23510 => "0000000000000000", 23511 => "0000000000000000", 23512 => "0000000000000000", 23513 => "0000000000000000", 23514 => "0000000000000000", 23515 => "0000000000000000", 23516 => "0000000000000000", 23517 => "0000000000000000", 23518 => "0000000000000000", 23519 => "0000000000000000", 23520 => "0000000000000000", 23521 => "0000000000000000", 23522 => "0000000000000000", 23523 => "0000000000000000", 23524 => "0000000000000000", 23525 => "0000000000000000", 23526 => "0000000000000000", 23527 => "0000000000000000", 23528 => "0000000000000000", 23529 => "0000000000000000", 23530 => "0000000000000000", 23531 => "0000000000000000", 23532 => "0000000000000000", 23533 => "0000000000000000", 23534 => "0000000000000000", 23535 => "0000000000000000", 23536 => "0000000000000000", 23537 => "0000000000000000", 23538 => "0000000000000000", 23539 => "0000000000000000", 23540 => "0000000000000000", 23541 => "0000000000000000", 23542 => "0000000000000000", 23543 => "0000000000000000", 23544 => "0000000000000000", 23545 => "0000000000000000", 23546 => "0000000000000000", 23547 => "0000000000000000", 23548 => "0000000000000000", 23549 => "0000000000000000", 23550 => "0000000000000000", 23551 => "0000000000000000", 23552 => "0000000000000000", 23553 => "0000000000000000", 23554 => "0000000000000000", 23555 => "0000000000000000", 23556 => "0000000000000000", 23557 => "0000000000000000", 23558 => "0000000000000000", 23559 => "0000000000000000", 23560 => "0000000000000000", 23561 => "0000000000000000", 23562 => "0000000000000000", 23563 => "0000000000000000", 23564 => "0000000000000000", 23565 => "0000000000000000", 23566 => "0000000000000000", 23567 => "0000000000000000", 23568 => "0000000000000000", 23569 => "0000000000000000", 23570 => "0000000000000000", 23571 => "0000000000000000", 23572 => "0000000000000000", 23573 => "0000000000000000", 23574 => "0000000000000000", 23575 => "0000000000000000", 23576 => "0000000000000000", 23577 => "0000000000000000", 23578 => "0000000000000000", 23579 => "0000000000000000", 23580 => "0000000000000000", 23581 => "0000000000000000", 23582 => "0000000000000000", 23583 => "0000000000000000", 23584 => "0000000000000000", 23585 => "0000000000000000", 23586 => "0000000000000000", 23587 => "0000000000000000", 23588 => "0000000000000000", 23589 => "0000000000000000", 23590 => "0000000000000000", 23591 => "0000000000000000", 23592 => "0000000000000000", 23593 => "0000000000000000", 23594 => "0000000000000000", 23595 => "0000000000000000", 23596 => "0000000000000000", 23597 => "0000000000000000", 23598 => "0000000000000000", 23599 => "0000000000000000", 23600 => "0000000000000000", 23601 => "0000000000000000", 23602 => "0000000000000000", 23603 => "0000000000000000", 23604 => "0000000000000000", 23605 => "0000000000000000", 23606 => "0000000000000000", 23607 => "0000000000000000", 23608 => "0000000000000000", 23609 => "0000000000000000", 23610 => "0000000000000000", 23611 => "0000000000000000", 23612 => "0000000000000000", 23613 => "0000000000000000", 23614 => "0000000000000000", 23615 => "0000000000000000", 23616 => "0000000000000000", 23617 => "0000000000000000", 23618 => "0000000000000000", 23619 => "0000000000000000", 23620 => "0000000000000000", 23621 => "0000000000000000", 23622 => "0000000000000000", 23623 => "0000000000000000", 23624 => "0000000000000000", 23625 => "0000000000000000", 23626 => "0000000000000000", 23627 => "0000000000000000", 23628 => "0000000000000000", 23629 => "0000000000000000", 23630 => "0000000000000000", 23631 => "0000000000000000", 23632 => "0000000000000000", 23633 => "0000000000000000", 23634 => "0000000000000000", 23635 => "0000000000000000", 23636 => "0000000000000000", 23637 => "0000000000000000", 23638 => "0000000000000000", 23639 => "0000000000000000", 23640 => "0000000000000000", 23641 => "0000000000000000", 23642 => "0000000000000000", 23643 => "0000000000000000", 23644 => "0000000000000000", 23645 => "0000000000000000", 23646 => "0000000000000000", 23647 => "0000000000000000", 23648 => "0000000000000000", 23649 => "0000000000000000", 23650 => "0000000000000000", 23651 => "0000000000000000", 23652 => "0000000000000000", 23653 => "0000000000000000", 23654 => "0000000000000000", 23655 => "0000000000000000", 23656 => "0000000000000000", 23657 => "0000000000000000", 23658 => "0000000000000000", 23659 => "0000000000000000", 23660 => "0000000000000000", 23661 => "0000000000000000", 23662 => "0000000000000000", 23663 => "0000000000000000", 23664 => "0000000000000000", 23665 => "0000000000000000", 23666 => "0000000000000000", 23667 => "0000000000000000", 23668 => "0000000000000000", 23669 => "0000000000000000", 23670 => "0000000000000000", 23671 => "0000000000000000", 23672 => "0000000000000000", 23673 => "0000000000000000", 23674 => "0000000000000000", 23675 => "0000000000000000", 23676 => "0000000000000000", 23677 => "0000000000000000", 23678 => "0000000000000000", 23679 => "0000000000000000", 23680 => "0000000000000000", 23681 => "0000000000000000", 23682 => "0000000000000000", 23683 => "0000000000000000", 23684 => "0000000000000000", 23685 => "0000000000000000", 23686 => "0000000000000000", 23687 => "0000000000000000", 23688 => "0000000000000000", 23689 => "0000000000000000", 23690 => "0000000000000000", 23691 => "0000000000000000", 23692 => "0000000000000000", 23693 => "0000000000000000", 23694 => "0000000000000000", 23695 => "0000000000000000", 23696 => "0000000000000000", 23697 => "0000000000000000", 23698 => "0000000000000000", 23699 => "0000000000000000", 23700 => "0000000000000000", 23701 => "0000000000000000", 23702 => "0000000000000000", 23703 => "0000000000000000", 23704 => "0000000000000000", 23705 => "0000000000000000", 23706 => "0000000000000000", 23707 => "0000000000000000", 23708 => "0000000000000000", 23709 => "0000000000000000", 23710 => "0000000000000000", 23711 => "0000000000000000", 23712 => "0000000000000000", 23713 => "0000000000000000", 23714 => "0000000000000000", 23715 => "0000000000000000", 23716 => "0000000000000000", 23717 => "0000000000000000", 23718 => "0000000000000000", 23719 => "0000000000000000", 23720 => "0000000000000000", 23721 => "0000000000000000", 23722 => "0000000000000000", 23723 => "0000000000000000", 23724 => "0000000000000000", 23725 => "0000000000000000", 23726 => "0000000000000000", 23727 => "0000000000000000", 23728 => "0000000000000000", 23729 => "0000000000000000", 23730 => "0000000000000000", 23731 => "0000000000000000", 23732 => "0000000000000000", 23733 => "0000000000000000", 23734 => "0000000000000000", 23735 => "0000000000000000", 23736 => "0000000000000000", 23737 => "0000000000000000", 23738 => "0000000000000000", 23739 => "0000000000000000", 23740 => "0000000000000000", 23741 => "0000000000000000", 23742 => "0000000000000000", 23743 => "0000000000000000", 23744 => "0000000000000000", 23745 => "0000000000000000", 23746 => "0000000000000000", 23747 => "0000000000000000", 23748 => "0000000000000000", 23749 => "0000000000000000", 23750 => "0000000000000000", 23751 => "0000000000000000", 23752 => "0000000000000000", 23753 => "0000000000000000", 23754 => "0000000000000000", 23755 => "0000000000000000", 23756 => "0000000000000000", 23757 => "0000000000000000", 23758 => "0000000000000000", 23759 => "0000000000000000", 23760 => "0000000000000000", 23761 => "0000000000000000", 23762 => "0000000000000000", 23763 => "0000000000000000", 23764 => "0000000000000000", 23765 => "0000000000000000", 23766 => "0000000000000000", 23767 => "0000000000000000", 23768 => "0000000000000000", 23769 => "0000000000000000", 23770 => "0000000000000000", 23771 => "0000000000000000", 23772 => "0000000000000000", 23773 => "0000000000000000", 23774 => "0000000000000000", 23775 => "0000000000000000", 23776 => "0000000000000000", 23777 => "0000000000000000", 23778 => "0000000000000000", 23779 => "0000000000000000", 23780 => "0000000000000000", 23781 => "0000000000000000", 23782 => "0000000000000000", 23783 => "0000000000000000", 23784 => "0000000000000000", 23785 => "0000000000000000", 23786 => "0000000000000000", 23787 => "0000000000000000", 23788 => "0000000000000000", 23789 => "0000000000000000", 23790 => "0000000000000000", 23791 => "0000000000000000", 23792 => "0000000000000000", 23793 => "0000000000000000", 23794 => "0000000000000000", 23795 => "0000000000000000", 23796 => "0000000000000000", 23797 => "0000000000000000", 23798 => "0000000000000000", 23799 => "0000000000000000", 23800 => "0000000000000000", 23801 => "0000000000000000", 23802 => "0000000000000000", 23803 => "0000000000000000", 23804 => "0000000000000000", 23805 => "0000000000000000", 23806 => "0000000000000000", 23807 => "0000000000000000", 23808 => "0000000000000000", 23809 => "0000000000000000", 23810 => "0000000000000000", 23811 => "0000000000000000", 23812 => "0000000000000000", 23813 => "0000000000000000", 23814 => "0000000000000000", 23815 => "0000000000000000", 23816 => "0000000000000000", 23817 => "0000000000000000", 23818 => "0000000000000000", 23819 => "0000000000000000", 23820 => "0000000000000000", 23821 => "0000000000000000", 23822 => "0000000000000000", 23823 => "0000000000000000", 23824 => "0000000000000000", 23825 => "0000000000000000", 23826 => "0000000000000000", 23827 => "0000000000000000", 23828 => "0000000000000000", 23829 => "0000000000000000", 23830 => "0000000000000000", 23831 => "0000000000000000", 23832 => "0000000000000000", 23833 => "0000000000000000", 23834 => "0000000000000000", 23835 => "0000000000000000", 23836 => "0000000000000000", 23837 => "0000000000000000", 23838 => "0000000000000000", 23839 => "0000000000000000", 23840 => "0000000000000000", 23841 => "0000000000000000", 23842 => "0000000000000000", 23843 => "0000000000000000", 23844 => "0000000000000000", 23845 => "0000000000000000", 23846 => "0000000000000000", 23847 => "0000000000000000", 23848 => "0000000000000000", 23849 => "0000000000000000", 23850 => "0000000000000000", 23851 => "0000000000000000", 23852 => "0000000000000000", 23853 => "0000000000000000", 23854 => "0000000000000000", 23855 => "0000000000000000", 23856 => "0000000000000000", 23857 => "0000000000000000", 23858 => "0000000000000000", 23859 => "0000000000000000", 23860 => "0000000000000000", 23861 => "0000000000000000", 23862 => "0000000000000000", 23863 => "0000000000000000", 23864 => "0000000000000000", 23865 => "0000000000000000", 23866 => "0000000000000000", 23867 => "0000000000000000", 23868 => "0000000000000000", 23869 => "0000000000000000", 23870 => "0000000000000000", 23871 => "0000000000000000", 23872 => "0000000000000000", 23873 => "0000000000000000", 23874 => "0000000000000000", 23875 => "0000000000000000", 23876 => "0000000000000000", 23877 => "0000000000000000", 23878 => "0000000000000000", 23879 => "0000000000000000", 23880 => "0000000000000000", 23881 => "0000000000000000", 23882 => "0000000000000000", 23883 => "0000000000000000", 23884 => "0000000000000000", 23885 => "0000000000000000", 23886 => "0000000000000000", 23887 => "0000000000000000", 23888 => "0000000000000000", 23889 => "0000000000000000", 23890 => "0000000000000000", 23891 => "0000000000000000", 23892 => "0000000000000000", 23893 => "0000000000000000", 23894 => "0000000000000000", 23895 => "0000000000000000", 23896 => "0000000000000000", 23897 => "0000000000000000", 23898 => "0000000000000000", 23899 => "0000000000000000", 23900 => "0000000000000000", 23901 => "0000000000000000", 23902 => "0000000000000000", 23903 => "0000000000000000", 23904 => "0000000000000000", 23905 => "0000000000000000", 23906 => "0000000000000000", 23907 => "0000000000000000", 23908 => "0000000000000000", 23909 => "0000000000000000", 23910 => "0000000000000000", 23911 => "0000000000000000", 23912 => "0000000000000000", 23913 => "0000000000000000", 23914 => "0000000000000000", 23915 => "0000000000000000", 23916 => "0000000000000000", 23917 => "0000000000000000", 23918 => "0000000000000000", 23919 => "0000000000000000", 23920 => "0000000000000000", 23921 => "0000000000000000", 23922 => "0000000000000000", 23923 => "0000000000000000", 23924 => "0000000000000000", 23925 => "0000000000000000", 23926 => "0000000000000000", 23927 => "0000000000000000", 23928 => "0000000000000000", 23929 => "0000000000000000", 23930 => "0000000000000000", 23931 => "0000000000000000", 23932 => "0000000000000000", 23933 => "0000000000000000", 23934 => "0000000000000000", 23935 => "0000000000000000", 23936 => "0000000000000000", 23937 => "0000000000000000", 23938 => "0000000000000000", 23939 => "0000000000000000", 23940 => "0000000000000000", 23941 => "0000000000000000", 23942 => "0000000000000000", 23943 => "0000000000000000", 23944 => "0000000000000000", 23945 => "0000000000000000", 23946 => "0000000000000000", 23947 => "0000000000000000", 23948 => "0000000000000000", 23949 => "0000000000000000", 23950 => "0000000000000000", 23951 => "0000000000000000", 23952 => "0000000000000000", 23953 => "0000000000000000", 23954 => "0000000000000000", 23955 => "0000000000000000", 23956 => "0000000000000000", 23957 => "0000000000000000", 23958 => "0000000000000000", 23959 => "0000000000000000", 23960 => "0000000000000000", 23961 => "0000000000000000", 23962 => "0000000000000000", 23963 => "0000000000000000", 23964 => "0000000000000000", 23965 => "0000000000000000", 23966 => "0000000000000000", 23967 => "0000000000000000", 23968 => "0000000000000000", 23969 => "0000000000000000", 23970 => "0000000000000000", 23971 => "0000000000000000", 23972 => "0000000000000000", 23973 => "0000000000000000", 23974 => "0000000000000000", 23975 => "0000000000000000", 23976 => "0000000000000000", 23977 => "0000000000000000", 23978 => "0000000000000000", 23979 => "0000000000000000", 23980 => "0000000000000000", 23981 => "0000000000000000", 23982 => "0000000000000000", 23983 => "0000000000000000", 23984 => "0000000000000000", 23985 => "0000000000000000", 23986 => "0000000000000000", 23987 => "0000000000000000", 23988 => "0000000000000000", 23989 => "0000000000000000", 23990 => "0000000000000000", 23991 => "0000000000000000", 23992 => "0000000000000000", 23993 => "0000000000000000", 23994 => "0000000000000000", 23995 => "0000000000000000", 23996 => "0000000000000000", 23997 => "0000000000000000", 23998 => "0000000000000000", 23999 => "0000000000000000", 24000 => "0000000000000000", 24001 => "0000000000000000", 24002 => "0000000000000000", 24003 => "0000000000000000", 24004 => "0000000000000000", 24005 => "0000000000000000", 24006 => "0000000000000000", 24007 => "0000000000000000", 24008 => "0000000000000000", 24009 => "0000000000000000", 24010 => "0000000000000000", 24011 => "0000000000000000", 24012 => "0000000000000000", 24013 => "0000000000000000", 24014 => "0000000000000000", 24015 => "0000000000000000", 24016 => "0000000000000000", 24017 => "0000000000000000", 24018 => "0000000000000000", 24019 => "0000000000000000", 24020 => "0000000000000000", 24021 => "0000000000000000", 24022 => "0000000000000000", 24023 => "0000000000000000", 24024 => "0000000000000000", 24025 => "0000000000000000", 24026 => "0000000000000000", 24027 => "0000000000000000", 24028 => "0000000000000000", 24029 => "0000000000000000", 24030 => "0000000000000000", 24031 => "0000000000000000", 24032 => "0000000000000000", 24033 => "0000000000000000", 24034 => "0000000000000000", 24035 => "0000000000000000", 24036 => "0000000000000000", 24037 => "0000000000000000", 24038 => "0000000000000000", 24039 => "0000000000000000", 24040 => "0000000000000000", 24041 => "0000000000000000", 24042 => "0000000000000000", 24043 => "0000000000000000", 24044 => "0000000000000000", 24045 => "0000000000000000", 24046 => "0000000000000000", 24047 => "0000000000000000", 24048 => "0000000000000000", 24049 => "0000000000000000", 24050 => "0000000000000000", 24051 => "0000000000000000", 24052 => "0000000000000000", 24053 => "0000000000000000", 24054 => "0000000000000000", 24055 => "0000000000000000", 24056 => "0000000000000000", 24057 => "0000000000000000", 24058 => "0000000000000000", 24059 => "0000000000000000", 24060 => "0000000000000000", 24061 => "0000000000000000", 24062 => "0000000000000000", 24063 => "0000000000000000", 24064 => "0000000000000000", 24065 => "0000000000000000", 24066 => "0000000000000000", 24067 => "0000000000000000", 24068 => "0000000000000000", 24069 => "0000000000000000", 24070 => "0000000000000000", 24071 => "0000000000000000", 24072 => "0000000000000000", 24073 => "0000000000000000", 24074 => "0000000000000000", 24075 => "0000000000000000", 24076 => "0000000000000000", 24077 => "0000000000000000", 24078 => "0000000000000000", 24079 => "0000000000000000", 24080 => "0000000000000000", 24081 => "0000000000000000", 24082 => "0000000000000000", 24083 => "0000000000000000", 24084 => "0000000000000000", 24085 => "0000000000000000", 24086 => "0000000000000000", 24087 => "0000000000000000", 24088 => "0000000000000000", 24089 => "0000000000000000", 24090 => "0000000000000000", 24091 => "0000000000000000", 24092 => "0000000000000000", 24093 => "0000000000000000", 24094 => "0000000000000000", 24095 => "0000000000000000", 24096 => "0000000000000000", 24097 => "0000000000000000", 24098 => "0000000000000000", 24099 => "0000000000000000", 24100 => "0000000000000000", 24101 => "0000000000000000", 24102 => "0000000000000000", 24103 => "0000000000000000", 24104 => "0000000000000000", 24105 => "0000000000000000", 24106 => "0000000000000000", 24107 => "0000000000000000", 24108 => "0000000000000000", 24109 => "0000000000000000", 24110 => "0000000000000000", 24111 => "0000000000000000", 24112 => "0000000000000000", 24113 => "0000000000000000", 24114 => "0000000000000000", 24115 => "0000000000000000", 24116 => "0000000000000000", 24117 => "0000000000000000", 24118 => "0000000000000000", 24119 => "0000000000000000", 24120 => "0000000000000000", 24121 => "0000000000000000", 24122 => "0000000000000000", 24123 => "0000000000000000", 24124 => "0000000000000000", 24125 => "0000000000000000", 24126 => "0000000000000000", 24127 => "0000000000000000", 24128 => "0000000000000000", 24129 => "0000000000000000", 24130 => "0000000000000000", 24131 => "0000000000000000", 24132 => "0000000000000000", 24133 => "0000000000000000", 24134 => "0000000000000000", 24135 => "0000000000000000", 24136 => "0000000000000000", 24137 => "0000000000000000", 24138 => "0000000000000000", 24139 => "0000000000000000", 24140 => "0000000000000000", 24141 => "0000000000000000", 24142 => "0000000000000000", 24143 => "0000000000000000", 24144 => "0000000000000000", 24145 => "0000000000000000", 24146 => "0000000000000000", 24147 => "0000000000000000", 24148 => "0000000000000000", 24149 => "0000000000000000", 24150 => "0000000000000000", 24151 => "0000000000000000", 24152 => "0000000000000000", 24153 => "0000000000000000", 24154 => "0000000000000000", 24155 => "0000000000000000", 24156 => "0000000000000000", 24157 => "0000000000000000", 24158 => "0000000000000000", 24159 => "0000000000000000", 24160 => "0000000000000000", 24161 => "0000000000000000", 24162 => "0000000000000000", 24163 => "0000000000000000", 24164 => "0000000000000000", 24165 => "0000000000000000", 24166 => "0000000000000000", 24167 => "0000000000000000", 24168 => "0000000000000000", 24169 => "0000000000000000", 24170 => "0000000000000000", 24171 => "0000000000000000", 24172 => "0000000000000000", 24173 => "0000000000000000", 24174 => "0000000000000000", 24175 => "0000000000000000", 24176 => "0000000000000000", 24177 => "0000000000000000", 24178 => "0000000000000000", 24179 => "0000000000000000", 24180 => "0000000000000000", 24181 => "0000000000000000", 24182 => "0000000000000000", 24183 => "0000000000000000", 24184 => "0000000000000000", 24185 => "0000000000000000", 24186 => "0000000000000000", 24187 => "0000000000000000", 24188 => "0000000000000000", 24189 => "0000000000000000", 24190 => "0000000000000000", 24191 => "0000000000000000", 24192 => "0000000000000000", 24193 => "0000000000000000", 24194 => "0000000000000000", 24195 => "0000000000000000", 24196 => "0000000000000000", 24197 => "0000000000000000", 24198 => "0000000000000000", 24199 => "0000000000000000", 24200 => "0000000000000000", 24201 => "0000000000000000", 24202 => "0000000000000000", 24203 => "0000000000000000", 24204 => "0000000000000000", 24205 => "0000000000000000", 24206 => "0000000000000000", 24207 => "0000000000000000", 24208 => "0000000000000000", 24209 => "0000000000000000", 24210 => "0000000000000000", 24211 => "0000000000000000", 24212 => "0000000000000000", 24213 => "0000000000000000", 24214 => "0000000000000000", 24215 => "0000000000000000", 24216 => "0000000000000000", 24217 => "0000000000000000", 24218 => "0000000000000000", 24219 => "0000000000000000", 24220 => "0000000000000000", 24221 => "0000000000000000", 24222 => "0000000000000000", 24223 => "0000000000000000", 24224 => "0000000000000000", 24225 => "0000000000000000", 24226 => "0000000000000000", 24227 => "0000000000000000", 24228 => "0000000000000000", 24229 => "0000000000000000", 24230 => "0000000000000000", 24231 => "0000000000000000", 24232 => "0000000000000000", 24233 => "0000000000000000", 24234 => "0000000000000000", 24235 => "0000000000000000", 24236 => "0000000000000000", 24237 => "0000000000000000", 24238 => "0000000000000000", 24239 => "0000000000000000", 24240 => "0000000000000000", 24241 => "0000000000000000", 24242 => "0000000000000000", 24243 => "0000000000000000", 24244 => "0000000000000000", 24245 => "0000000000000000", 24246 => "0000000000000000", 24247 => "0000000000000000", 24248 => "0000000000000000", 24249 => "0000000000000000", 24250 => "0000000000000000", 24251 => "0000000000000000", 24252 => "0000000000000000", 24253 => "0000000000000000", 24254 => "0000000000000000", 24255 => "0000000000000000", 24256 => "0000000000000000", 24257 => "0000000000000000", 24258 => "0000000000000000", 24259 => "0000000000000000", 24260 => "0000000000000000", 24261 => "0000000000000000", 24262 => "0000000000000000", 24263 => "0000000000000000", 24264 => "0000000000000000", 24265 => "0000000000000000", 24266 => "0000000000000000", 24267 => "0000000000000000", 24268 => "0000000000000000", 24269 => "0000000000000000", 24270 => "0000000000000000", 24271 => "0000000000000000", 24272 => "0000000000000000", 24273 => "0000000000000000", 24274 => "0000000000000000", 24275 => "0000000000000000", 24276 => "0000000000000000", 24277 => "0000000000000000", 24278 => "0000000000000000", 24279 => "0000000000000000", 24280 => "0000000000000000", 24281 => "0000000000000000", 24282 => "0000000000000000", 24283 => "0000000000000000", 24284 => "0000000000000000", 24285 => "0000000000000000", 24286 => "0000000000000000", 24287 => "0000000000000000", 24288 => "0000000000000000", 24289 => "0000000000000000", 24290 => "0000000000000000", 24291 => "0000000000000000", 24292 => "0000000000000000", 24293 => "0000000000000000", 24294 => "0000000000000000", 24295 => "0000000000000000", 24296 => "0000000000000000", 24297 => "0000000000000000", 24298 => "0000000000000000", 24299 => "0000000000000000", 24300 => "0000000000000000", 24301 => "0000000000000000", 24302 => "0000000000000000", 24303 => "0000000000000000", 24304 => "0000000000000000", 24305 => "0000000000000000", 24306 => "0000000000000000", 24307 => "0000000000000000", 24308 => "0000000000000000", 24309 => "0000000000000000", 24310 => "0000000000000000", 24311 => "0000000000000000", 24312 => "0000000000000000", 24313 => "0000000000000000", 24314 => "0000000000000000", 24315 => "0000000000000000", 24316 => "0000000000000000", 24317 => "0000000000000000", 24318 => "0000000000000000", 24319 => "0000000000000000", 24320 => "0000000000000000", 24321 => "0000000000000000", 24322 => "0000000000000000", 24323 => "0000000000000000", 24324 => "0000000000000000", 24325 => "0000000000000000", 24326 => "0000000000000000", 24327 => "0000000000000000", 24328 => "0000000000000000", 24329 => "0000000000000000", 24330 => "0000000000000000", 24331 => "0000000000000000", 24332 => "0000000000000000", 24333 => "0000000000000000", 24334 => "0000000000000000", 24335 => "0000000000000000", 24336 => "0000000000000000", 24337 => "0000000000000000", 24338 => "0000000000000000", 24339 => "0000000000000000", 24340 => "0000000000000000", 24341 => "0000000000000000", 24342 => "0000000000000000", 24343 => "0000000000000000", 24344 => "0000000000000000", 24345 => "0000000000000000", 24346 => "0000000000000000", 24347 => "0000000000000000", 24348 => "0000000000000000", 24349 => "0000000000000000", 24350 => "0000000000000000", 24351 => "0000000000000000", 24352 => "0000000000000000", 24353 => "0000000000000000", 24354 => "0000000000000000", 24355 => "0000000000000000", 24356 => "0000000000000000", 24357 => "0000000000000000", 24358 => "0000000000000000", 24359 => "0000000000000000", 24360 => "0000000000000000", 24361 => "0000000000000000", 24362 => "0000000000000000", 24363 => "0000000000000000", 24364 => "0000000000000000", 24365 => "0000000000000000", 24366 => "0000000000000000", 24367 => "0000000000000000", 24368 => "0000000000000000", 24369 => "0000000000000000", 24370 => "0000000000000000", 24371 => "0000000000000000", 24372 => "0000000000000000", 24373 => "0000000000000000", 24374 => "0000000000000000", 24375 => "0000000000000000", 24376 => "0000000000000000", 24377 => "0000000000000000", 24378 => "0000000000000000", 24379 => "0000000000000000", 24380 => "0000000000000000", 24381 => "0000000000000000", 24382 => "0000000000000000", 24383 => "0000000000000000", 24384 => "0000000000000000", 24385 => "0000000000000000", 24386 => "0000000000000000", 24387 => "0000000000000000", 24388 => "0000000000000000", 24389 => "0000000000000000", 24390 => "0000000000000000", 24391 => "0000000000000000", 24392 => "0000000000000000", 24393 => "0000000000000000", 24394 => "0000000000000000", 24395 => "0000000000000000", 24396 => "0000000000000000", 24397 => "0000000000000000", 24398 => "0000000000000000", 24399 => "0000000000000000", 24400 => "0000000000000000", 24401 => "0000000000000000", 24402 => "0000000000000000", 24403 => "0000000000000000", 24404 => "0000000000000000", 24405 => "0000000000000000", 24406 => "0000000000000000", 24407 => "0000000000000000", 24408 => "0000000000000000", 24409 => "0000000000000000", 24410 => "0000000000000000", 24411 => "0000000000000000", 24412 => "0000000000000000", 24413 => "0000000000000000", 24414 => "0000000000000000", 24415 => "0000000000000000", 24416 => "0000000000000000", 24417 => "0000000000000000", 24418 => "0000000000000000", 24419 => "0000000000000000", 24420 => "0000000000000000", 24421 => "0000000000000000", 24422 => "0000000000000000", 24423 => "0000000000000000", 24424 => "0000000000000000", 24425 => "0000000000000000", 24426 => "0000000000000000", 24427 => "0000000000000000", 24428 => "0000000000000000", 24429 => "0000000000000000", 24430 => "0000000000000000", 24431 => "0000000000000000", 24432 => "0000000000000000", 24433 => "0000000000000000", 24434 => "0000000000000000", 24435 => "0000000000000000", 24436 => "0000000000000000", 24437 => "0000000000000000", 24438 => "0000000000000000", 24439 => "0000000000000000", 24440 => "0000000000000000", 24441 => "0000000000000000", 24442 => "0000000000000000", 24443 => "0000000000000000", 24444 => "0000000000000000", 24445 => "0000000000000000", 24446 => "0000000000000000", 24447 => "0000000000000000", 24448 => "0000000000000000", 24449 => "0000000000000000", 24450 => "0000000000000000", 24451 => "0000000000000000", 24452 => "0000000000000000", 24453 => "0000000000000000", 24454 => "0000000000000000", 24455 => "0000000000000000", 24456 => "0000000000000000", 24457 => "0000000000000000", 24458 => "0000000000000000", 24459 => "0000000000000000", 24460 => "0000000000000000", 24461 => "0000000000000000", 24462 => "0000000000000000", 24463 => "0000000000000000", 24464 => "0000000000000000", 24465 => "0000000000000000", 24466 => "0000000000000000", 24467 => "0000000000000000", 24468 => "0000000000000000", 24469 => "0000000000000000", 24470 => "0000000000000000", 24471 => "0000000000000000", 24472 => "0000000000000000", 24473 => "0000000000000000", 24474 => "0000000000000000", 24475 => "0000000000000000", 24476 => "0000000000000000", 24477 => "0000000000000000", 24478 => "0000000000000000", 24479 => "0000000000000000", 24480 => "0000000000000000", 24481 => "0000000000000000", 24482 => "0000000000000000", 24483 => "0000000000000000", 24484 => "0000000000000000", 24485 => "0000000000000000", 24486 => "0000000000000000", 24487 => "0000000000000000", 24488 => "0000000000000000", 24489 => "0000000000000000", 24490 => "0000000000000000", 24491 => "0000000000000000", 24492 => "0000000000000000", 24493 => "0000000000000000", 24494 => "0000000000000000", 24495 => "0000000000000000", 24496 => "0000000000000000", 24497 => "0000000000000000", 24498 => "0000000000000000", 24499 => "0000000000000000", 24500 => "0000000000000000", 24501 => "0000000000000000", 24502 => "0000000000000000", 24503 => "0000000000000000", 24504 => "0000000000000000", 24505 => "0000000000000000", 24506 => "0000000000000000", 24507 => "0000000000000000", 24508 => "0000000000000000", 24509 => "0000000000000000", 24510 => "0000000000000000", 24511 => "0000000000000000", 24512 => "0000000000000000", 24513 => "0000000000000000", 24514 => "0000000000000000", 24515 => "0000000000000000", 24516 => "0000000000000000", 24517 => "0000000000000000", 24518 => "0000000000000000", 24519 => "0000000000000000", 24520 => "0000000000000000", 24521 => "0000000000000000", 24522 => "0000000000000000", 24523 => "0000000000000000", 24524 => "0000000000000000", 24525 => "0000000000000000", 24526 => "0000000000000000", 24527 => "0000000000000000", 24528 => "0000000000000000", 24529 => "0000000000000000", 24530 => "0000000000000000", 24531 => "0000000000000000", 24532 => "0000000000000000", 24533 => "0000000000000000", 24534 => "0000000000000000", 24535 => "0000000000000000", 24536 => "0000000000000000", 24537 => "0000000000000000", 24538 => "0000000000000000", 24539 => "0000000000000000", 24540 => "0000000000000000", 24541 => "0000000000000000", 24542 => "0000000000000000", 24543 => "0000000000000000", 24544 => "0000000000000000", 24545 => "0000000000000000", 24546 => "0000000000000000", 24547 => "0000000000000000", 24548 => "0000000000000000", 24549 => "0000000000000000", 24550 => "0000000000000000", 24551 => "0000000000000000", 24552 => "0000000000000000", 24553 => "0000000000000000", 24554 => "0000000000000000", 24555 => "0000000000000000", 24556 => "0000000000000000", 24557 => "0000000000000000", 24558 => "0000000000000000", 24559 => "0000000000000000", 24560 => "0000000000000000", 24561 => "0000000000000000", 24562 => "0000000000000000", 24563 => "0000000000000000", 24564 => "0000000000000000", 24565 => "0000000000000000", 24566 => "0000000000000000", 24567 => "0000000000000000", 24568 => "0000000000000000", 24569 => "0000000000000000", 24570 => "0000000000000000", 24571 => "0000000000000000", 24572 => "0000000000000000", 24573 => "0000000000000000", 24574 => "0000000000000000", 24575 => "0000000000000000", 24576 => "0000000000000000", 24577 => "0000000000000000", 24578 => "0000000000000000", 24579 => "0000000000000000", 24580 => "0000000000000000", 24581 => "0000000000000000", 24582 => "0000000000000000", 24583 => "0000000000000000", 24584 => "0000000000000000", 24585 => "0000000000000000", 24586 => "0000000000000000", 24587 => "0000000000000000", 24588 => "0000000000000000", 24589 => "0000000000000000", 24590 => "0000000000000000", 24591 => "0000000000000000", 24592 => "0000000000000000", 24593 => "0000000000000000", 24594 => "0000000000000000", 24595 => "0000000000000000", 24596 => "0000000000000000", 24597 => "0000000000000000", 24598 => "0000000000000000", 24599 => "0000000000000000", 24600 => "0000000000000000", 24601 => "0000000000000000", 24602 => "0000000000000000", 24603 => "0000000000000000", 24604 => "0000000000000000", 24605 => "0000000000000000", 24606 => "0000000000000000", 24607 => "0000000000000000", 24608 => "0000000000000000", 24609 => "0000000000000000", 24610 => "0000000000000000", 24611 => "0000000000000000", 24612 => "0000000000000000", 24613 => "0000000000000000", 24614 => "0000000000000000", 24615 => "0000000000000000", 24616 => "0000000000000000", 24617 => "0000000000000000", 24618 => "0000000000000000", 24619 => "0000000000000000", 24620 => "0000000000000000", 24621 => "0000000000000000", 24622 => "0000000000000000", 24623 => "0000000000000000", 24624 => "0000000000000000", 24625 => "0000000000000000", 24626 => "0000000000000000", 24627 => "0000000000000000", 24628 => "0000000000000000", 24629 => "0000000000000000", 24630 => "0000000000000000", 24631 => "0000000000000000", 24632 => "0000000000000000", 24633 => "0000000000000000", 24634 => "0000000000000000", 24635 => "0000000000000000", 24636 => "0000000000000000", 24637 => "0000000000000000", 24638 => "0000000000000000", 24639 => "0000000000000000", 24640 => "0000000000000000", 24641 => "0000000000000000", 24642 => "0000000000000000", 24643 => "0000000000000000", 24644 => "0000000000000000", 24645 => "0000000000000000", 24646 => "0000000000000000", 24647 => "0000000000000000", 24648 => "0000000000000000", 24649 => "0000000000000000", 24650 => "0000000000000000", 24651 => "0000000000000000", 24652 => "0000000000000000", 24653 => "0000000000000000", 24654 => "0000000000000000", 24655 => "0000000000000000", 24656 => "0000000000000000", 24657 => "0000000000000000", 24658 => "0000000000000000", 24659 => "0000000000000000", 24660 => "0000000000000000", 24661 => "0000000000000000", 24662 => "0000000000000000", 24663 => "0000000000000000", 24664 => "0000000000000000", 24665 => "0000000000000000", 24666 => "0000000000000000", 24667 => "0000000000000000", 24668 => "0000000000000000", 24669 => "0000000000000000", 24670 => "0000000000000000", 24671 => "0000000000000000", 24672 => "0000000000000000", 24673 => "0000000000000000", 24674 => "0000000000000000", 24675 => "0000000000000000", 24676 => "0000000000000000", 24677 => "0000000000000000", 24678 => "0000000000000000", 24679 => "0000000000000000", 24680 => "0000000000000000", 24681 => "0000000000000000", 24682 => "0000000000000000", 24683 => "0000000000000000", 24684 => "0000000000000000", 24685 => "0000000000000000", 24686 => "0000000000000000", 24687 => "0000000000000000", 24688 => "0000000000000000", 24689 => "0000000000000000", 24690 => "0000000000000000", 24691 => "0000000000000000", 24692 => "0000000000000000", 24693 => "0000000000000000", 24694 => "0000000000000000", 24695 => "0000000000000000", 24696 => "0000000000000000", 24697 => "0000000000000000", 24698 => "0000000000000000", 24699 => "0000000000000000", 24700 => "0000000000000000", 24701 => "0000000000000000", 24702 => "0000000000000000", 24703 => "0000000000000000", 24704 => "0000000000000000", 24705 => "0000000000000000", 24706 => "0000000000000000", 24707 => "0000000000000000", 24708 => "0000000000000000", 24709 => "0000000000000000", 24710 => "0000000000000000", 24711 => "0000000000000000", 24712 => "0000000000000000", 24713 => "0000000000000000", 24714 => "0000000000000000", 24715 => "0000000000000000", 24716 => "0000000000000000", 24717 => "0000000000000000", 24718 => "0000000000000000", 24719 => "0000000000000000", 24720 => "0000000000000000", 24721 => "0000000000000000", 24722 => "0000000000000000", 24723 => "0000000000000000", 24724 => "0000000000000000", 24725 => "0000000000000000", 24726 => "0000000000000000", 24727 => "0000000000000000", 24728 => "0000000000000000", 24729 => "0000000000000000", 24730 => "0000000000000000", 24731 => "0000000000000000", 24732 => "0000000000000000", 24733 => "0000000000000000", 24734 => "0000000000000000", 24735 => "0000000000000000", 24736 => "0000000000000000", 24737 => "0000000000000000", 24738 => "0000000000000000", 24739 => "0000000000000000", 24740 => "0000000000000000", 24741 => "0000000000000000", 24742 => "0000000000000000", 24743 => "0000000000000000", 24744 => "0000000000000000", 24745 => "0000000000000000", 24746 => "0000000000000000", 24747 => "0000000000000000", 24748 => "0000000000000000", 24749 => "0000000000000000", 24750 => "0000000000000000", 24751 => "0000000000000000", 24752 => "0000000000000000", 24753 => "0000000000000000", 24754 => "0000000000000000", 24755 => "0000000000000000", 24756 => "0000000000000000", 24757 => "0000000000000000", 24758 => "0000000000000000", 24759 => "0000000000000000", 24760 => "0000000000000000", 24761 => "0000000000000000", 24762 => "0000000000000000", 24763 => "0000000000000000", 24764 => "0000000000000000", 24765 => "0000000000000000", 24766 => "0000000000000000", 24767 => "0000000000000000", 24768 => "0000000000000000", 24769 => "0000000000000000", 24770 => "0000000000000000", 24771 => "0000000000000000", 24772 => "0000000000000000", 24773 => "0000000000000000", 24774 => "0000000000000000", 24775 => "0000000000000000", 24776 => "0000000000000000", 24777 => "0000000000000000", 24778 => "0000000000000000", 24779 => "0000000000000000", 24780 => "0000000000000000", 24781 => "0000000000000000", 24782 => "0000000000000000", 24783 => "0000000000000000", 24784 => "0000000000000000", 24785 => "0000000000000000", 24786 => "0000000000000000", 24787 => "0000000000000000", 24788 => "0000000000000000", 24789 => "0000000000000000", 24790 => "0000000000000000", 24791 => "0000000000000000", 24792 => "0000000000000000", 24793 => "0000000000000000", 24794 => "0000000000000000", 24795 => "0000000000000000", 24796 => "0000000000000000", 24797 => "0000000000000000", 24798 => "0000000000000000", 24799 => "0000000000000000", 24800 => "0000000000000000", 24801 => "0000000000000000", 24802 => "0000000000000000", 24803 => "0000000000000000", 24804 => "0000000000000000", 24805 => "0000000000000000", 24806 => "0000000000000000", 24807 => "0000000000000000", 24808 => "0000000000000000", 24809 => "0000000000000000", 24810 => "0000000000000000", 24811 => "0000000000000000", 24812 => "0000000000000000", 24813 => "0000000000000000", 24814 => "0000000000000000", 24815 => "0000000000000000", 24816 => "0000000000000000", 24817 => "0000000000000000", 24818 => "0000000000000000", 24819 => "0000000000000000", 24820 => "0000000000000000", 24821 => "0000000000000000", 24822 => "0000000000000000", 24823 => "0000000000000000", 24824 => "0000000000000000", 24825 => "0000000000000000", 24826 => "0000000000000000", 24827 => "0000000000000000", 24828 => "0000000000000000", 24829 => "0000000000000000", 24830 => "0000000000000000", 24831 => "0000000000000000", 24832 => "0000000000000000", 24833 => "0000000000000000", 24834 => "0000000000000000", 24835 => "0000000000000000", 24836 => "0000000000000000", 24837 => "0000000000000000", 24838 => "0000000000000000", 24839 => "0000000000000000", 24840 => "0000000000000000", 24841 => "0000000000000000", 24842 => "0000000000000000", 24843 => "0000000000000000", 24844 => "0000000000000000", 24845 => "0000000000000000", 24846 => "0000000000000000", 24847 => "0000000000000000", 24848 => "0000000000000000", 24849 => "0000000000000000", 24850 => "0000000000000000", 24851 => "0000000000000000", 24852 => "0000000000000000", 24853 => "0000000000000000", 24854 => "0000000000000000", 24855 => "0000000000000000", 24856 => "0000000000000000", 24857 => "0000000000000000", 24858 => "0000000000000000", 24859 => "0000000000000000", 24860 => "0000000000000000", 24861 => "0000000000000000", 24862 => "0000000000000000", 24863 => "0000000000000000", 24864 => "0000000000000000", 24865 => "0000000000000000", 24866 => "0000000000000000", 24867 => "0000000000000000", 24868 => "0000000000000000", 24869 => "0000000000000000", 24870 => "0000000000000000", 24871 => "0000000000000000", 24872 => "0000000000000000", 24873 => "0000000000000000", 24874 => "0000000000000000", 24875 => "0000000000000000", 24876 => "0000000000000000", 24877 => "0000000000000000", 24878 => "0000000000000000", 24879 => "0000000000000000", 24880 => "0000000000000000", 24881 => "0000000000000000", 24882 => "0000000000000000", 24883 => "0000000000000000", 24884 => "0000000000000000", 24885 => "0000000000000000", 24886 => "0000000000000000", 24887 => "0000000000000000", 24888 => "0000000000000000", 24889 => "0000000000000000", 24890 => "0000000000000000", 24891 => "0000000000000000", 24892 => "0000000000000000", 24893 => "0000000000000000", 24894 => "0000000000000000", 24895 => "0000000000000000", 24896 => "0000000000000000", 24897 => "0000000000000000", 24898 => "0000000000000000", 24899 => "0000000000000000", 24900 => "0000000000000000", 24901 => "0000000000000000", 24902 => "0000000000000000", 24903 => "0000000000000000", 24904 => "0000000000000000", 24905 => "0000000000000000", 24906 => "0000000000000000", 24907 => "0000000000000000", 24908 => "0000000000000000", 24909 => "0000000000000000", 24910 => "0000000000000000", 24911 => "0000000000000000", 24912 => "0000000000000000", 24913 => "0000000000000000", 24914 => "0000000000000000", 24915 => "0000000000000000", 24916 => "0000000000000000", 24917 => "0000000000000000", 24918 => "0000000000000000", 24919 => "0000000000000000", 24920 => "0000000000000000", 24921 => "0000000000000000", 24922 => "0000000000000000", 24923 => "0000000000000000", 24924 => "0000000000000000", 24925 => "0000000000000000", 24926 => "0000000000000000", 24927 => "0000000000000000", 24928 => "0000000000000000", 24929 => "0000000000000000", 24930 => "0000000000000000", 24931 => "0000000000000000", 24932 => "0000000000000000", 24933 => "0000000000000000", 24934 => "0000000000000000", 24935 => "0000000000000000", 24936 => "0000000000000000", 24937 => "0000000000000000", 24938 => "0000000000000000", 24939 => "0000000000000000", 24940 => "0000000000000000", 24941 => "0000000000000000", 24942 => "0000000000000000", 24943 => "0000000000000000", 24944 => "0000000000000000", 24945 => "0000000000000000", 24946 => "0000000000000000", 24947 => "0000000000000000", 24948 => "0000000000000000", 24949 => "0000000000000000", 24950 => "0000000000000000", 24951 => "0000000000000000", 24952 => "0000000000000000", 24953 => "0000000000000000", 24954 => "0000000000000000", 24955 => "0000000000000000", 24956 => "0000000000000000", 24957 => "0000000000000000", 24958 => "0000000000000000", 24959 => "0000000000000000", 24960 => "0000000000000000", 24961 => "0000000000000000", 24962 => "0000000000000000", 24963 => "0000000000000000", 24964 => "0000000000000000", 24965 => "0000000000000000", 24966 => "0000000000000000", 24967 => "0000000000000000", 24968 => "0000000000000000", 24969 => "0000000000000000", 24970 => "0000000000000000", 24971 => "0000000000000000", 24972 => "0000000000000000", 24973 => "0000000000000000", 24974 => "0000000000000000", 24975 => "0000000000000000", 24976 => "0000000000000000", 24977 => "0000000000000000", 24978 => "0000000000000000", 24979 => "0000000000000000", 24980 => "0000000000000000", 24981 => "0000000000000000", 24982 => "0000000000000000", 24983 => "0000000000000000", 24984 => "0000000000000000", 24985 => "0000000000000000", 24986 => "0000000000000000", 24987 => "0000000000000000", 24988 => "0000000000000000", 24989 => "0000000000000000", 24990 => "0000000000000000", 24991 => "0000000000000000", 24992 => "0000000000000000", 24993 => "0000000000000000", 24994 => "0000000000000000", 24995 => "0000000000000000", 24996 => "0000000000000000", 24997 => "0000000000000000", 24998 => "0000000000000000", 24999 => "0000000000000000", 25000 => "0000000000000000", 25001 => "0000000000000000", 25002 => "0000000000000000", 25003 => "0000000000000000", 25004 => "0000000000000000", 25005 => "0000000000000000", 25006 => "0000000000000000", 25007 => "0000000000000000", 25008 => "0000000000000000", 25009 => "0000000000000000", 25010 => "0000000000000000", 25011 => "0000000000000000", 25012 => "0000000000000000", 25013 => "0000000000000000", 25014 => "0000000000000000", 25015 => "0000000000000000", 25016 => "0000000000000000", 25017 => "0000000000000000", 25018 => "0000000000000000", 25019 => "0000000000000000", 25020 => "0000000000000000", 25021 => "0000000000000000", 25022 => "0000000000000000", 25023 => "0000000000000000", 25024 => "0000000000000000", 25025 => "0000000000000000", 25026 => "0000000000000000", 25027 => "0000000000000000", 25028 => "0000000000000000", 25029 => "0000000000000000", 25030 => "0000000000000000", 25031 => "0000000000000000", 25032 => "0000000000000000", 25033 => "0000000000000000", 25034 => "0000000000000000", 25035 => "0000000000000000", 25036 => "0000000000000000", 25037 => "0000000000000000", 25038 => "0000000000000000", 25039 => "0000000000000000", 25040 => "0000000000000000", 25041 => "0000000000000000", 25042 => "0000000000000000", 25043 => "0000000000000000", 25044 => "0000000000000000", 25045 => "0000000000000000", 25046 => "0000000000000000", 25047 => "0000000000000000", 25048 => "0000000000000000", 25049 => "0000000000000000", 25050 => "0000000000000000", 25051 => "0000000000000000", 25052 => "0000000000000000", 25053 => "0000000000000000", 25054 => "0000000000000000", 25055 => "0000000000000000", 25056 => "0000000000000000", 25057 => "0000000000000000", 25058 => "0000000000000000", 25059 => "0000000000000000", 25060 => "0000000000000000", 25061 => "0000000000000000", 25062 => "0000000000000000", 25063 => "0000000000000000", 25064 => "0000000000000000", 25065 => "0000000000000000", 25066 => "0000000000000000", 25067 => "0000000000000000", 25068 => "0000000000000000", 25069 => "0000000000000000", 25070 => "0000000000000000", 25071 => "0000000000000000", 25072 => "0000000000000000", 25073 => "0000000000000000", 25074 => "0000000000000000", 25075 => "0000000000000000", 25076 => "0000000000000000", 25077 => "0000000000000000", 25078 => "0000000000000000", 25079 => "0000000000000000", 25080 => "0000000000000000", 25081 => "0000000000000000", 25082 => "0000000000000000", 25083 => "0000000000000000", 25084 => "0000000000000000", 25085 => "0000000000000000", 25086 => "0000000000000000", 25087 => "0000000000000000", 25088 => "0000000000000000", 25089 => "0000000000000000", 25090 => "0000000000000000", 25091 => "0000000000000000", 25092 => "0000000000000000", 25093 => "0000000000000000", 25094 => "0000000000000000", 25095 => "0000000000000000", 25096 => "0000000000000000", 25097 => "0000000000000000", 25098 => "0000000000000000", 25099 => "0000000000000000", 25100 => "0000000000000000", 25101 => "0000000000000000", 25102 => "0000000000000000", 25103 => "0000000000000000", 25104 => "0000000000000000", 25105 => "0000000000000000", 25106 => "0000000000000000", 25107 => "0000000000000000", 25108 => "0000000000000000", 25109 => "0000000000000000", 25110 => "0000000000000000", 25111 => "0000000000000000", 25112 => "0000000000000000", 25113 => "0000000000000000", 25114 => "0000000000000000", 25115 => "0000000000000000", 25116 => "0000000000000000", 25117 => "0000000000000000", 25118 => "0000000000000000", 25119 => "0000000000000000", 25120 => "0000000000000000", 25121 => "0000000000000000", 25122 => "0000000000000000", 25123 => "0000000000000000", 25124 => "0000000000000000", 25125 => "0000000000000000", 25126 => "0000000000000000", 25127 => "0000000000000000", 25128 => "0000000000000000", 25129 => "0000000000000000", 25130 => "0000000000000000", 25131 => "0000000000000000", 25132 => "0000000000000000", 25133 => "0000000000000000", 25134 => "0000000000000000", 25135 => "0000000000000000", 25136 => "0000000000000000", 25137 => "0000000000000000", 25138 => "0000000000000000", 25139 => "0000000000000000", 25140 => "0000000000000000", 25141 => "0000000000000000", 25142 => "0000000000000000", 25143 => "0000000000000000", 25144 => "0000000000000000", 25145 => "0000000000000000", 25146 => "0000000000000000", 25147 => "0000000000000000", 25148 => "0000000000000000", 25149 => "0000000000000000", 25150 => "0000000000000000", 25151 => "0000000000000000", 25152 => "0000000000000000", 25153 => "0000000000000000", 25154 => "0000000000000000", 25155 => "0000000000000000", 25156 => "0000000000000000", 25157 => "0000000000000000", 25158 => "0000000000000000", 25159 => "0000000000000000", 25160 => "0000000000000000", 25161 => "0000000000000000", 25162 => "0000000000000000", 25163 => "0000000000000000", 25164 => "0000000000000000", 25165 => "0000000000000000", 25166 => "0000000000000000", 25167 => "0000000000000000", 25168 => "0000000000000000", 25169 => "0000000000000000", 25170 => "0000000000000000", 25171 => "0000000000000000", 25172 => "0000000000000000", 25173 => "0000000000000000", 25174 => "0000000000000000", 25175 => "0000000000000000", 25176 => "0000000000000000", 25177 => "0000000000000000", 25178 => "0000000000000000", 25179 => "0000000000000000", 25180 => "0000000000000000", 25181 => "0000000000000000", 25182 => "0000000000000000", 25183 => "0000000000000000", 25184 => "0000000000000000", 25185 => "0000000000000000", 25186 => "0000000000000000", 25187 => "0000000000000000", 25188 => "0000000000000000", 25189 => "0000000000000000", 25190 => "0000000000000000", 25191 => "0000000000000000", 25192 => "0000000000000000", 25193 => "0000000000000000", 25194 => "0000000000000000", 25195 => "0000000000000000", 25196 => "0000000000000000", 25197 => "0000000000000000", 25198 => "0000000000000000", 25199 => "0000000000000000", 25200 => "0000000000000000", 25201 => "0000000000000000", 25202 => "0000000000000000", 25203 => "0000000000000000", 25204 => "0000000000000000", 25205 => "0000000000000000", 25206 => "0000000000000000", 25207 => "0000000000000000", 25208 => "0000000000000000", 25209 => "0000000000000000", 25210 => "0000000000000000", 25211 => "0000000000000000", 25212 => "0000000000000000", 25213 => "0000000000000000", 25214 => "0000000000000000", 25215 => "0000000000000000", 25216 => "0000000000000000", 25217 => "0000000000000000", 25218 => "0000000000000000", 25219 => "0000000000000000", 25220 => "0000000000000000", 25221 => "0000000000000000", 25222 => "0000000000000000", 25223 => "0000000000000000", 25224 => "0000000000000000", 25225 => "0000000000000000", 25226 => "0000000000000000", 25227 => "0000000000000000", 25228 => "0000000000000000", 25229 => "0000000000000000", 25230 => "0000000000000000", 25231 => "0000000000000000", 25232 => "0000000000000000", 25233 => "0000000000000000", 25234 => "0000000000000000", 25235 => "0000000000000000", 25236 => "0000000000000000", 25237 => "0000000000000000", 25238 => "0000000000000000", 25239 => "0000000000000000", 25240 => "0000000000000000", 25241 => "0000000000000000", 25242 => "0000000000000000", 25243 => "0000000000000000", 25244 => "0000000000000000", 25245 => "0000000000000000", 25246 => "0000000000000000", 25247 => "0000000000000000", 25248 => "0000000000000000", 25249 => "0000000000000000", 25250 => "0000000000000000", 25251 => "0000000000000000", 25252 => "0000000000000000", 25253 => "0000000000000000", 25254 => "0000000000000000", 25255 => "0000000000000000", 25256 => "0000000000000000", 25257 => "0000000000000000", 25258 => "0000000000000000", 25259 => "0000000000000000", 25260 => "0000000000000000", 25261 => "0000000000000000", 25262 => "0000000000000000", 25263 => "0000000000000000", 25264 => "0000000000000000", 25265 => "0000000000000000", 25266 => "0000000000000000", 25267 => "0000000000000000", 25268 => "0000000000000000", 25269 => "0000000000000000", 25270 => "0000000000000000", 25271 => "0000000000000000", 25272 => "0000000000000000", 25273 => "0000000000000000", 25274 => "0000000000000000", 25275 => "0000000000000000", 25276 => "0000000000000000", 25277 => "0000000000000000", 25278 => "0000000000000000", 25279 => "0000000000000000", 25280 => "0000000000000000", 25281 => "0000000000000000", 25282 => "0000000000000000", 25283 => "0000000000000000", 25284 => "0000000000000000", 25285 => "0000000000000000", 25286 => "0000000000000000", 25287 => "0000000000000000", 25288 => "0000000000000000", 25289 => "0000000000000000", 25290 => "0000000000000000", 25291 => "0000000000000000", 25292 => "0000000000000000", 25293 => "0000000000000000", 25294 => "0000000000000000", 25295 => "0000000000000000", 25296 => "0000000000000000", 25297 => "0000000000000000", 25298 => "0000000000000000", 25299 => "0000000000000000", 25300 => "0000000000000000", 25301 => "0000000000000000", 25302 => "0000000000000000", 25303 => "0000000000000000", 25304 => "0000000000000000", 25305 => "0000000000000000", 25306 => "0000000000000000", 25307 => "0000000000000000", 25308 => "0000000000000000", 25309 => "0000000000000000", 25310 => "0000000000000000", 25311 => "0000000000000000", 25312 => "0000000000000000", 25313 => "0000000000000000", 25314 => "0000000000000000", 25315 => "0000000000000000", 25316 => "0000000000000000", 25317 => "0000000000000000", 25318 => "0000000000000000", 25319 => "0000000000000000", 25320 => "0000000000000000", 25321 => "0000000000000000", 25322 => "0000000000000000", 25323 => "0000000000000000", 25324 => "0000000000000000", 25325 => "0000000000000000", 25326 => "0000000000000000", 25327 => "0000000000000000", 25328 => "0000000000000000", 25329 => "0000000000000000", 25330 => "0000000000000000", 25331 => "0000000000000000", 25332 => "0000000000000000", 25333 => "0000000000000000", 25334 => "0000000000000000", 25335 => "0000000000000000", 25336 => "0000000000000000", 25337 => "0000000000000000", 25338 => "0000000000000000", 25339 => "0000000000000000", 25340 => "0000000000000000", 25341 => "0000000000000000", 25342 => "0000000000000000", 25343 => "0000000000000000", 25344 => "0000000000000000", 25345 => "0000000000000000", 25346 => "0000000000000000", 25347 => "0000000000000000", 25348 => "0000000000000000", 25349 => "0000000000000000", 25350 => "0000000000000000", 25351 => "0000000000000000", 25352 => "0000000000000000", 25353 => "0000000000000000", 25354 => "0000000000000000", 25355 => "0000000000000000", 25356 => "0000000000000000", 25357 => "0000000000000000", 25358 => "0000000000000000", 25359 => "0000000000000000", 25360 => "0000000000000000", 25361 => "0000000000000000", 25362 => "0000000000000000", 25363 => "0000000000000000", 25364 => "0000000000000000", 25365 => "0000000000000000", 25366 => "0000000000000000", 25367 => "0000000000000000", 25368 => "0000000000000000", 25369 => "0000000000000000", 25370 => "0000000000000000", 25371 => "0000000000000000", 25372 => "0000000000000000", 25373 => "0000000000000000", 25374 => "0000000000000000", 25375 => "0000000000000000", 25376 => "0000000000000000", 25377 => "0000000000000000", 25378 => "0000000000000000", 25379 => "0000000000000000", 25380 => "0000000000000000", 25381 => "0000000000000000", 25382 => "0000000000000000", 25383 => "0000000000000000", 25384 => "0000000000000000", 25385 => "0000000000000000", 25386 => "0000000000000000", 25387 => "0000000000000000", 25388 => "0000000000000000", 25389 => "0000000000000000", 25390 => "0000000000000000", 25391 => "0000000000000000", 25392 => "0000000000000000", 25393 => "0000000000000000", 25394 => "0000000000000000", 25395 => "0000000000000000", 25396 => "0000000000000000", 25397 => "0000000000000000", 25398 => "0000000000000000", 25399 => "0000000000000000", 25400 => "0000000000000000", 25401 => "0000000000000000", 25402 => "0000000000000000", 25403 => "0000000000000000", 25404 => "0000000000000000", 25405 => "0000000000000000", 25406 => "0000000000000000", 25407 => "0000000000000000", 25408 => "0000000000000000", 25409 => "0000000000000000", 25410 => "0000000000000000", 25411 => "0000000000000000", 25412 => "0000000000000000", 25413 => "0000000000000000", 25414 => "0000000000000000", 25415 => "0000000000000000", 25416 => "0000000000000000", 25417 => "0000000000000000", 25418 => "0000000000000000", 25419 => "0000000000000000", 25420 => "0000000000000000", 25421 => "0000000000000000", 25422 => "0000000000000000", 25423 => "0000000000000000", 25424 => "0000000000000000", 25425 => "0000000000000000", 25426 => "0000000000000000", 25427 => "0000000000000000", 25428 => "0000000000000000", 25429 => "0000000000000000", 25430 => "0000000000000000", 25431 => "0000000000000000", 25432 => "0000000000000000", 25433 => "0000000000000000", 25434 => "0000000000000000", 25435 => "0000000000000000", 25436 => "0000000000000000", 25437 => "0000000000000000", 25438 => "0000000000000000", 25439 => "0000000000000000", 25440 => "0000000000000000", 25441 => "0000000000000000", 25442 => "0000000000000000", 25443 => "0000000000000000", 25444 => "0000000000000000", 25445 => "0000000000000000", 25446 => "0000000000000000", 25447 => "0000000000000000", 25448 => "0000000000000000", 25449 => "0000000000000000", 25450 => "0000000000000000", 25451 => "0000000000000000", 25452 => "0000000000000000", 25453 => "0000000000000000", 25454 => "0000000000000000", 25455 => "0000000000000000", 25456 => "0000000000000000", 25457 => "0000000000000000", 25458 => "0000000000000000", 25459 => "0000000000000000", 25460 => "0000000000000000", 25461 => "0000000000000000", 25462 => "0000000000000000", 25463 => "0000000000000000", 25464 => "0000000000000000", 25465 => "0000000000000000", 25466 => "0000000000000000", 25467 => "0000000000000000", 25468 => "0000000000000000", 25469 => "0000000000000000", 25470 => "0000000000000000", 25471 => "0000000000000000", 25472 => "0000000000000000", 25473 => "0000000000000000", 25474 => "0000000000000000", 25475 => "0000000000000000", 25476 => "0000000000000000", 25477 => "0000000000000000", 25478 => "0000000000000000", 25479 => "0000000000000000", 25480 => "0000000000000000", 25481 => "0000000000000000", 25482 => "0000000000000000", 25483 => "0000000000000000", 25484 => "0000000000000000", 25485 => "0000000000000000", 25486 => "0000000000000000", 25487 => "0000000000000000", 25488 => "0000000000000000", 25489 => "0000000000000000", 25490 => "0000000000000000", 25491 => "0000000000000000", 25492 => "0000000000000000", 25493 => "0000000000000000", 25494 => "0000000000000000", 25495 => "0000000000000000", 25496 => "0000000000000000", 25497 => "0000000000000000", 25498 => "0000000000000000", 25499 => "0000000000000000", 25500 => "0000000000000000", 25501 => "0000000000000000", 25502 => "0000000000000000", 25503 => "0000000000000000", 25504 => "0000000000000000", 25505 => "0000000000000000", 25506 => "0000000000000000", 25507 => "0000000000000000", 25508 => "0000000000000000", 25509 => "0000000000000000", 25510 => "0000000000000000", 25511 => "0000000000000000", 25512 => "0000000000000000", 25513 => "0000000000000000", 25514 => "0000000000000000", 25515 => "0000000000000000", 25516 => "0000000000000000", 25517 => "0000000000000000", 25518 => "0000000000000000", 25519 => "0000000000000000", 25520 => "0000000000000000", 25521 => "0000000000000000", 25522 => "0000000000000000", 25523 => "0000000000000000", 25524 => "0000000000000000", 25525 => "0000000000000000", 25526 => "0000000000000000", 25527 => "0000000000000000", 25528 => "0000000000000000", 25529 => "0000000000000000", 25530 => "0000000000000000", 25531 => "0000000000000000", 25532 => "0000000000000000", 25533 => "0000000000000000", 25534 => "0000000000000000", 25535 => "0000000000000000", 25536 => "0000000000000000", 25537 => "0000000000000000", 25538 => "0000000000000000", 25539 => "0000000000000000", 25540 => "0000000000000000", 25541 => "0000000000000000", 25542 => "0000000000000000", 25543 => "0000000000000000", 25544 => "0000000000000000", 25545 => "0000000000000000", 25546 => "0000000000000000", 25547 => "0000000000000000", 25548 => "0000000000000000", 25549 => "0000000000000000", 25550 => "0000000000000000", 25551 => "0000000000000000", 25552 => "0000000000000000", 25553 => "0000000000000000", 25554 => "0000000000000000", 25555 => "0000000000000000", 25556 => "0000000000000000", 25557 => "0000000000000000", 25558 => "0000000000000000", 25559 => "0000000000000000", 25560 => "0000000000000000", 25561 => "0000000000000000", 25562 => "0000000000000000", 25563 => "0000000000000000", 25564 => "0000000000000000", 25565 => "0000000000000000", 25566 => "0000000000000000", 25567 => "0000000000000000", 25568 => "0000000000000000", 25569 => "0000000000000000", 25570 => "0000000000000000", 25571 => "0000000000000000", 25572 => "0000000000000000", 25573 => "0000000000000000", 25574 => "0000000000000000", 25575 => "0000000000000000", 25576 => "0000000000000000", 25577 => "0000000000000000", 25578 => "0000000000000000", 25579 => "0000000000000000", 25580 => "0000000000000000", 25581 => "0000000000000000", 25582 => "0000000000000000", 25583 => "0000000000000000", 25584 => "0000000000000000", 25585 => "0000000000000000", 25586 => "0000000000000000", 25587 => "0000000000000000", 25588 => "0000000000000000", 25589 => "0000000000000000", 25590 => "0000000000000000", 25591 => "0000000000000000", 25592 => "0000000000000000", 25593 => "0000000000000000", 25594 => "0000000000000000", 25595 => "0000000000000000", 25596 => "0000000000000000", 25597 => "0000000000000000", 25598 => "0000000000000000", 25599 => "0000000000000000", 25600 => "0000000000000000", 25601 => "0000000000000000", 25602 => "0000000000000000", 25603 => "0000000000000000", 25604 => "0000000000000000", 25605 => "0000000000000000", 25606 => "0000000000000000", 25607 => "0000000000000000", 25608 => "0000000000000000", 25609 => "0000000000000000", 25610 => "0000000000000000", 25611 => "0000000000000000", 25612 => "0000000000000000", 25613 => "0000000000000000", 25614 => "0000000000000000", 25615 => "0000000000000000", 25616 => "0000000000000000", 25617 => "0000000000000000", 25618 => "0000000000000000", 25619 => "0000000000000000", 25620 => "0000000000000000", 25621 => "0000000000000000", 25622 => "0000000000000000", 25623 => "0000000000000000", 25624 => "0000000000000000", 25625 => "0000000000000000", 25626 => "0000000000000000", 25627 => "0000000000000000", 25628 => "0000000000000000", 25629 => "0000000000000000", 25630 => "0000000000000000", 25631 => "0000000000000000", 25632 => "0000000000000000", 25633 => "0000000000000000", 25634 => "0000000000000000", 25635 => "0000000000000000", 25636 => "0000000000000000", 25637 => "0000000000000000", 25638 => "0000000000000000", 25639 => "0000000000000000", 25640 => "0000000000000000", 25641 => "0000000000000000", 25642 => "0000000000000000", 25643 => "0000000000000000", 25644 => "0000000000000000", 25645 => "0000000000000000", 25646 => "0000000000000000", 25647 => "0000000000000000", 25648 => "0000000000000000", 25649 => "0000000000000000", 25650 => "0000000000000000", 25651 => "0000000000000000", 25652 => "0000000000000000", 25653 => "0000000000000000", 25654 => "0000000000000000", 25655 => "0000000000000000", 25656 => "0000000000000000", 25657 => "0000000000000000", 25658 => "0000000000000000", 25659 => "0000000000000000", 25660 => "0000000000000000", 25661 => "0000000000000000", 25662 => "0000000000000000", 25663 => "0000000000000000", 25664 => "0000000000000000", 25665 => "0000000000000000", 25666 => "0000000000000000", 25667 => "0000000000000000", 25668 => "0000000000000000", 25669 => "0000000000000000", 25670 => "0000000000000000", 25671 => "0000000000000000", 25672 => "0000000000000000", 25673 => "0000000000000000", 25674 => "0000000000000000", 25675 => "0000000000000000", 25676 => "0000000000000000", 25677 => "0000000000000000", 25678 => "0000000000000000", 25679 => "0000000000000000", 25680 => "0000000000000000", 25681 => "0000000000000000", 25682 => "0000000000000000", 25683 => "0000000000000000", 25684 => "0000000000000000", 25685 => "0000000000000000", 25686 => "0000000000000000", 25687 => "0000000000000000", 25688 => "0000000000000000", 25689 => "0000000000000000", 25690 => "0000000000000000", 25691 => "0000000000000000", 25692 => "0000000000000000", 25693 => "0000000000000000", 25694 => "0000000000000000", 25695 => "0000000000000000", 25696 => "0000000000000000", 25697 => "0000000000000000", 25698 => "0000000000000000", 25699 => "0000000000000000", 25700 => "0000000000000000", 25701 => "0000000000000000", 25702 => "0000000000000000", 25703 => "0000000000000000", 25704 => "0000000000000000", 25705 => "0000000000000000", 25706 => "0000000000000000", 25707 => "0000000000000000", 25708 => "0000000000000000", 25709 => "0000000000000000", 25710 => "0000000000000000", 25711 => "0000000000000000", 25712 => "0000000000000000", 25713 => "0000000000000000", 25714 => "0000000000000000", 25715 => "0000000000000000", 25716 => "0000000000000000", 25717 => "0000000000000000", 25718 => "0000000000000000", 25719 => "0000000000000000", 25720 => "0000000000000000", 25721 => "0000000000000000", 25722 => "0000000000000000", 25723 => "0000000000000000", 25724 => "0000000000000000", 25725 => "0000000000000000", 25726 => "0000000000000000", 25727 => "0000000000000000", 25728 => "0000000000000000", 25729 => "0000000000000000", 25730 => "0000000000000000", 25731 => "0000000000000000", 25732 => "0000000000000000", 25733 => "0000000000000000", 25734 => "0000000000000000", 25735 => "0000000000000000", 25736 => "0000000000000000", 25737 => "0000000000000000", 25738 => "0000000000000000", 25739 => "0000000000000000", 25740 => "0000000000000000", 25741 => "0000000000000000", 25742 => "0000000000000000", 25743 => "0000000000000000", 25744 => "0000000000000000", 25745 => "0000000000000000", 25746 => "0000000000000000", 25747 => "0000000000000000", 25748 => "0000000000000000", 25749 => "0000000000000000", 25750 => "0000000000000000", 25751 => "0000000000000000", 25752 => "0000000000000000", 25753 => "0000000000000000", 25754 => "0000000000000000", 25755 => "0000000000000000", 25756 => "0000000000000000", 25757 => "0000000000000000", 25758 => "0000000000000000", 25759 => "0000000000000000", 25760 => "0000000000000000", 25761 => "0000000000000000", 25762 => "0000000000000000", 25763 => "0000000000000000", 25764 => "0000000000000000", 25765 => "0000000000000000", 25766 => "0000000000000000", 25767 => "0000000000000000", 25768 => "0000000000000000", 25769 => "0000000000000000", 25770 => "0000000000000000", 25771 => "0000000000000000", 25772 => "0000000000000000", 25773 => "0000000000000000", 25774 => "0000000000000000", 25775 => "0000000000000000", 25776 => "0000000000000000", 25777 => "0000000000000000", 25778 => "0000000000000000", 25779 => "0000000000000000", 25780 => "0000000000000000", 25781 => "0000000000000000", 25782 => "0000000000000000", 25783 => "0000000000000000", 25784 => "0000000000000000", 25785 => "0000000000000000", 25786 => "0000000000000000", 25787 => "0000000000000000", 25788 => "0000000000000000", 25789 => "0000000000000000", 25790 => "0000000000000000", 25791 => "0000000000000000", 25792 => "0000000000000000", 25793 => "0000000000000000", 25794 => "0000000000000000", 25795 => "0000000000000000", 25796 => "0000000000000000", 25797 => "0000000000000000", 25798 => "0000000000000000", 25799 => "0000000000000000", 25800 => "0000000000000000", 25801 => "0000000000000000", 25802 => "0000000000000000", 25803 => "0000000000000000", 25804 => "0000000000000000", 25805 => "0000000000000000", 25806 => "0000000000000000", 25807 => "0000000000000000", 25808 => "0000000000000000", 25809 => "0000000000000000", 25810 => "0000000000000000", 25811 => "0000000000000000", 25812 => "0000000000000000", 25813 => "0000000000000000", 25814 => "0000000000000000", 25815 => "0000000000000000", 25816 => "0000000000000000", 25817 => "0000000000000000", 25818 => "0000000000000000", 25819 => "0000000000000000", 25820 => "0000000000000000", 25821 => "0000000000000000", 25822 => "0000000000000000", 25823 => "0000000000000000", 25824 => "0000000000000000", 25825 => "0000000000000000", 25826 => "0000000000000000", 25827 => "0000000000000000", 25828 => "0000000000000000", 25829 => "0000000000000000", 25830 => "0000000000000000", 25831 => "0000000000000000", 25832 => "0000000000000000", 25833 => "0000000000000000", 25834 => "0000000000000000", 25835 => "0000000000000000", 25836 => "0000000000000000", 25837 => "0000000000000000", 25838 => "0000000000000000", 25839 => "0000000000000000", 25840 => "0000000000000000", 25841 => "0000000000000000", 25842 => "0000000000000000", 25843 => "0000000000000000", 25844 => "0000000000000000", 25845 => "0000000000000000", 25846 => "0000000000000000", 25847 => "0000000000000000", 25848 => "0000000000000000", 25849 => "0000000000000000", 25850 => "0000000000000000", 25851 => "0000000000000000", 25852 => "0000000000000000", 25853 => "0000000000000000", 25854 => "0000000000000000", 25855 => "0000000000000000", 25856 => "0000000000000000", 25857 => "0000000000000000", 25858 => "0000000000000000", 25859 => "0000000000000000", 25860 => "0000000000000000", 25861 => "0000000000000000", 25862 => "0000000000000000", 25863 => "0000000000000000", 25864 => "0000000000000000", 25865 => "0000000000000000", 25866 => "0000000000000000", 25867 => "0000000000000000", 25868 => "0000000000000000", 25869 => "0000000000000000", 25870 => "0000000000000000", 25871 => "0000000000000000", 25872 => "0000000000000000", 25873 => "0000000000000000", 25874 => "0000000000000000", 25875 => "0000000000000000", 25876 => "0000000000000000", 25877 => "0000000000000000", 25878 => "0000000000000000", 25879 => "0000000000000000", 25880 => "0000000000000000", 25881 => "0000000000000000", 25882 => "0000000000000000", 25883 => "0000000000000000", 25884 => "0000000000000000", 25885 => "0000000000000000", 25886 => "0000000000000000", 25887 => "0000000000000000", 25888 => "0000000000000000", 25889 => "0000000000000000", 25890 => "0000000000000000", 25891 => "0000000000000000", 25892 => "0000000000000000", 25893 => "0000000000000000", 25894 => "0000000000000000", 25895 => "0000000000000000", 25896 => "0000000000000000", 25897 => "0000000000000000", 25898 => "0000000000000000", 25899 => "0000000000000000", 25900 => "0000000000000000", 25901 => "0000000000000000", 25902 => "0000000000000000", 25903 => "0000000000000000", 25904 => "0000000000000000", 25905 => "0000000000000000", 25906 => "0000000000000000", 25907 => "0000000000000000", 25908 => "0000000000000000", 25909 => "0000000000000000", 25910 => "0000000000000000", 25911 => "0000000000000000", 25912 => "0000000000000000", 25913 => "0000000000000000", 25914 => "0000000000000000", 25915 => "0000000000000000", 25916 => "0000000000000000", 25917 => "0000000000000000", 25918 => "0000000000000000", 25919 => "0000000000000000", 25920 => "0000000000000000", 25921 => "0000000000000000", 25922 => "0000000000000000", 25923 => "0000000000000000", 25924 => "0000000000000000", 25925 => "0000000000000000", 25926 => "0000000000000000", 25927 => "0000000000000000", 25928 => "0000000000000000", 25929 => "0000000000000000", 25930 => "0000000000000000", 25931 => "0000000000000000", 25932 => "0000000000000000", 25933 => "0000000000000000", 25934 => "0000000000000000", 25935 => "0000000000000000", 25936 => "0000000000000000", 25937 => "0000000000000000", 25938 => "0000000000000000", 25939 => "0000000000000000", 25940 => "0000000000000000", 25941 => "0000000000000000", 25942 => "0000000000000000", 25943 => "0000000000000000", 25944 => "0000000000000000", 25945 => "0000000000000000", 25946 => "0000000000000000", 25947 => "0000000000000000", 25948 => "0000000000000000", 25949 => "0000000000000000", 25950 => "0000000000000000", 25951 => "0000000000000000", 25952 => "0000000000000000", 25953 => "0000000000000000", 25954 => "0000000000000000", 25955 => "0000000000000000", 25956 => "0000000000000000", 25957 => "0000000000000000", 25958 => "0000000000000000", 25959 => "0000000000000000", 25960 => "0000000000000000", 25961 => "0000000000000000", 25962 => "0000000000000000", 25963 => "0000000000000000", 25964 => "0000000000000000", 25965 => "0000000000000000", 25966 => "0000000000000000", 25967 => "0000000000000000", 25968 => "0000000000000000", 25969 => "0000000000000000", 25970 => "0000000000000000", 25971 => "0000000000000000", 25972 => "0000000000000000", 25973 => "0000000000000000", 25974 => "0000000000000000", 25975 => "0000000000000000", 25976 => "0000000000000000", 25977 => "0000000000000000", 25978 => "0000000000000000", 25979 => "0000000000000000", 25980 => "0000000000000000", 25981 => "0000000000000000", 25982 => "0000000000000000", 25983 => "0000000000000000", 25984 => "0000000000000000", 25985 => "0000000000000000", 25986 => "0000000000000000", 25987 => "0000000000000000", 25988 => "0000000000000000", 25989 => "0000000000000000", 25990 => "0000000000000000", 25991 => "0000000000000000", 25992 => "0000000000000000", 25993 => "0000000000000000", 25994 => "0000000000000000", 25995 => "0000000000000000", 25996 => "0000000000000000", 25997 => "0000000000000000", 25998 => "0000000000000000", 25999 => "0000000000000000", 26000 => "0000000000000000", 26001 => "0000000000000000", 26002 => "0000000000000000", 26003 => "0000000000000000", 26004 => "0000000000000000", 26005 => "0000000000000000", 26006 => "0000000000000000", 26007 => "0000000000000000", 26008 => "0000000000000000", 26009 => "0000000000000000", 26010 => "0000000000000000", 26011 => "0000000000000000", 26012 => "0000000000000000", 26013 => "0000000000000000", 26014 => "0000000000000000", 26015 => "0000000000000000", 26016 => "0000000000000000", 26017 => "0000000000000000", 26018 => "0000000000000000", 26019 => "0000000000000000", 26020 => "0000000000000000", 26021 => "0000000000000000", 26022 => "0000000000000000", 26023 => "0000000000000000", 26024 => "0000000000000000", 26025 => "0000000000000000", 26026 => "0000000000000000", 26027 => "0000000000000000", 26028 => "0000000000000000", 26029 => "0000000000000000", 26030 => "0000000000000000", 26031 => "0000000000000000", 26032 => "0000000000000000", 26033 => "0000000000000000", 26034 => "0000000000000000", 26035 => "0000000000000000", 26036 => "0000000000000000", 26037 => "0000000000000000", 26038 => "0000000000000000", 26039 => "0000000000000000", 26040 => "0000000000000000", 26041 => "0000000000000000", 26042 => "0000000000000000", 26043 => "0000000000000000", 26044 => "0000000000000000", 26045 => "0000000000000000", 26046 => "0000000000000000", 26047 => "0000000000000000", 26048 => "0000000000000000", 26049 => "0000000000000000", 26050 => "0000000000000000", 26051 => "0000000000000000", 26052 => "0000000000000000", 26053 => "0000000000000000", 26054 => "0000000000000000", 26055 => "0000000000000000", 26056 => "0000000000000000", 26057 => "0000000000000000", 26058 => "0000000000000000", 26059 => "0000000000000000", 26060 => "0000000000000000", 26061 => "0000000000000000", 26062 => "0000000000000000", 26063 => "0000000000000000", 26064 => "0000000000000000", 26065 => "0000000000000000", 26066 => "0000000000000000", 26067 => "0000000000000000", 26068 => "0000000000000000", 26069 => "0000000000000000", 26070 => "0000000000000000", 26071 => "0000000000000000", 26072 => "0000000000000000", 26073 => "0000000000000000", 26074 => "0000000000000000", 26075 => "0000000000000000", 26076 => "0000000000000000", 26077 => "0000000000000000", 26078 => "0000000000000000", 26079 => "0000000000000000", 26080 => "0000000000000000", 26081 => "0000000000000000", 26082 => "0000000000000000", 26083 => "0000000000000000", 26084 => "0000000000000000", 26085 => "0000000000000000", 26086 => "0000000000000000", 26087 => "0000000000000000", 26088 => "0000000000000000", 26089 => "0000000000000000", 26090 => "0000000000000000", 26091 => "0000000000000000", 26092 => "0000000000000000", 26093 => "0000000000000000", 26094 => "0000000000000000", 26095 => "0000000000000000", 26096 => "0000000000000000", 26097 => "0000000000000000", 26098 => "0000000000000000", 26099 => "0000000000000000", 26100 => "0000000000000000", 26101 => "0000000000000000", 26102 => "0000000000000000", 26103 => "0000000000000000", 26104 => "0000000000000000", 26105 => "0000000000000000", 26106 => "0000000000000000", 26107 => "0000000000000000", 26108 => "0000000000000000", 26109 => "0000000000000000", 26110 => "0000000000000000", 26111 => "0000000000000000", 26112 => "0000000000000000", 26113 => "0000000000000000", 26114 => "0000000000000000", 26115 => "0000000000000000", 26116 => "0000000000000000", 26117 => "0000000000000000", 26118 => "0000000000000000", 26119 => "0000000000000000", 26120 => "0000000000000000", 26121 => "0000000000000000", 26122 => "0000000000000000", 26123 => "0000000000000000", 26124 => "0000000000000000", 26125 => "0000000000000000", 26126 => "0000000000000000", 26127 => "0000000000000000", 26128 => "0000000000000000", 26129 => "0000000000000000", 26130 => "0000000000000000", 26131 => "0000000000000000", 26132 => "0000000000000000", 26133 => "0000000000000000", 26134 => "0000000000000000", 26135 => "0000000000000000", 26136 => "0000000000000000", 26137 => "0000000000000000", 26138 => "0000000000000000", 26139 => "0000000000000000", 26140 => "0000000000000000", 26141 => "0000000000000000", 26142 => "0000000000000000", 26143 => "0000000000000000", 26144 => "0000000000000000", 26145 => "0000000000000000", 26146 => "0000000000000000", 26147 => "0000000000000000", 26148 => "0000000000000000", 26149 => "0000000000000000", 26150 => "0000000000000000", 26151 => "0000000000000000", 26152 => "0000000000000000", 26153 => "0000000000000000", 26154 => "0000000000000000", 26155 => "0000000000000000", 26156 => "0000000000000000", 26157 => "0000000000000000", 26158 => "0000000000000000", 26159 => "0000000000000000", 26160 => "0000000000000000", 26161 => "0000000000000000", 26162 => "0000000000000000", 26163 => "0000000000000000", 26164 => "0000000000000000", 26165 => "0000000000000000", 26166 => "0000000000000000", 26167 => "0000000000000000", 26168 => "0000000000000000", 26169 => "0000000000000000", 26170 => "0000000000000000", 26171 => "0000000000000000", 26172 => "0000000000000000", 26173 => "0000000000000000", 26174 => "0000000000000000", 26175 => "0000000000000000", 26176 => "0000000000000000", 26177 => "0000000000000000", 26178 => "0000000000000000", 26179 => "0000000000000000", 26180 => "0000000000000000", 26181 => "0000000000000000", 26182 => "0000000000000000", 26183 => "0000000000000000", 26184 => "0000000000000000", 26185 => "0000000000000000", 26186 => "0000000000000000", 26187 => "0000000000000000", 26188 => "0000000000000000", 26189 => "0000000000000000", 26190 => "0000000000000000", 26191 => "0000000000000000", 26192 => "0000000000000000", 26193 => "0000000000000000", 26194 => "0000000000000000", 26195 => "0000000000000000", 26196 => "0000000000000000", 26197 => "0000000000000000", 26198 => "0000000000000000", 26199 => "0000000000000000", 26200 => "0000000000000000", 26201 => "0000000000000000", 26202 => "0000000000000000", 26203 => "0000000000000000", 26204 => "0000000000000000", 26205 => "0000000000000000", 26206 => "0000000000000000", 26207 => "0000000000000000", 26208 => "0000000000000000", 26209 => "0000000000000000", 26210 => "0000000000000000", 26211 => "0000000000000000", 26212 => "0000000000000000", 26213 => "0000000000000000", 26214 => "0000000000000000", 26215 => "0000000000000000", 26216 => "0000000000000000", 26217 => "0000000000000000", 26218 => "0000000000000000", 26219 => "0000000000000000", 26220 => "0000000000000000", 26221 => "0000000000000000", 26222 => "0000000000000000", 26223 => "0000000000000000", 26224 => "0000000000000000", 26225 => "0000000000000000", 26226 => "0000000000000000", 26227 => "0000000000000000", 26228 => "0000000000000000", 26229 => "0000000000000000", 26230 => "0000000000000000", 26231 => "0000000000000000", 26232 => "0000000000000000", 26233 => "0000000000000000", 26234 => "0000000000000000", 26235 => "0000000000000000", 26236 => "0000000000000000", 26237 => "0000000000000000", 26238 => "0000000000000000", 26239 => "0000000000000000", 26240 => "0000000000000000", 26241 => "0000000000000000", 26242 => "0000000000000000", 26243 => "0000000000000000", 26244 => "0000000000000000", 26245 => "0000000000000000", 26246 => "0000000000000000", 26247 => "0000000000000000", 26248 => "0000000000000000", 26249 => "0000000000000000", 26250 => "0000000000000000", 26251 => "0000000000000000", 26252 => "0000000000000000", 26253 => "0000000000000000", 26254 => "0000000000000000", 26255 => "0000000000000000", 26256 => "0000000000000000", 26257 => "0000000000000000", 26258 => "0000000000000000", 26259 => "0000000000000000", 26260 => "0000000000000000", 26261 => "0000000000000000", 26262 => "0000000000000000", 26263 => "0000000000000000", 26264 => "0000000000000000", 26265 => "0000000000000000", 26266 => "0000000000000000", 26267 => "0000000000000000", 26268 => "0000000000000000", 26269 => "0000000000000000", 26270 => "0000000000000000", 26271 => "0000000000000000", 26272 => "0000000000000000", 26273 => "0000000000000000", 26274 => "0000000000000000", 26275 => "0000000000000000", 26276 => "0000000000000000", 26277 => "0000000000000000", 26278 => "0000000000000000", 26279 => "0000000000000000", 26280 => "0000000000000000", 26281 => "0000000000000000", 26282 => "0000000000000000", 26283 => "0000000000000000", 26284 => "0000000000000000", 26285 => "0000000000000000", 26286 => "0000000000000000", 26287 => "0000000000000000", 26288 => "0000000000000000", 26289 => "0000000000000000", 26290 => "0000000000000000", 26291 => "0000000000000000", 26292 => "0000000000000000", 26293 => "0000000000000000", 26294 => "0000000000000000", 26295 => "0000000000000000", 26296 => "0000000000000000", 26297 => "0000000000000000", 26298 => "0000000000000000", 26299 => "0000000000000000", 26300 => "0000000000000000", 26301 => "0000000000000000", 26302 => "0000000000000000", 26303 => "0000000000000000", 26304 => "0000000000000000", 26305 => "0000000000000000", 26306 => "0000000000000000", 26307 => "0000000000000000", 26308 => "0000000000000000", 26309 => "0000000000000000", 26310 => "0000000000000000", 26311 => "0000000000000000", 26312 => "0000000000000000", 26313 => "0000000000000000", 26314 => "0000000000000000", 26315 => "0000000000000000", 26316 => "0000000000000000", 26317 => "0000000000000000", 26318 => "0000000000000000", 26319 => "0000000000000000", 26320 => "0000000000000000", 26321 => "0000000000000000", 26322 => "0000000000000000", 26323 => "0000000000000000", 26324 => "0000000000000000", 26325 => "0000000000000000", 26326 => "0000000000000000", 26327 => "0000000000000000", 26328 => "0000000000000000", 26329 => "0000000000000000", 26330 => "0000000000000000", 26331 => "0000000000000000", 26332 => "0000000000000000", 26333 => "0000000000000000", 26334 => "0000000000000000", 26335 => "0000000000000000", 26336 => "0000000000000000", 26337 => "0000000000000000", 26338 => "0000000000000000", 26339 => "0000000000000000", 26340 => "0000000000000000", 26341 => "0000000000000000", 26342 => "0000000000000000", 26343 => "0000000000000000", 26344 => "0000000000000000", 26345 => "0000000000000000", 26346 => "0000000000000000", 26347 => "0000000000000000", 26348 => "0000000000000000", 26349 => "0000000000000000", 26350 => "0000000000000000", 26351 => "0000000000000000", 26352 => "0000000000000000", 26353 => "0000000000000000", 26354 => "0000000000000000", 26355 => "0000000000000000", 26356 => "0000000000000000", 26357 => "0000000000000000", 26358 => "0000000000000000", 26359 => "0000000000000000", 26360 => "0000000000000000", 26361 => "0000000000000000", 26362 => "0000000000000000", 26363 => "0000000000000000", 26364 => "0000000000000000", 26365 => "0000000000000000", 26366 => "0000000000000000", 26367 => "0000000000000000", 26368 => "0000000000000000", 26369 => "0000000000000000", 26370 => "0000000000000000", 26371 => "0000000000000000", 26372 => "0000000000000000", 26373 => "0000000000000000", 26374 => "0000000000000000", 26375 => "0000000000000000", 26376 => "0000000000000000", 26377 => "0000000000000000", 26378 => "0000000000000000", 26379 => "0000000000000000", 26380 => "0000000000000000", 26381 => "0000000000000000", 26382 => "0000000000000000", 26383 => "0000000000000000", 26384 => "0000000000000000", 26385 => "0000000000000000", 26386 => "0000000000000000", 26387 => "0000000000000000", 26388 => "0000000000000000", 26389 => "0000000000000000", 26390 => "0000000000000000", 26391 => "0000000000000000", 26392 => "0000000000000000", 26393 => "0000000000000000", 26394 => "0000000000000000", 26395 => "0000000000000000", 26396 => "0000000000000000", 26397 => "0000000000000000", 26398 => "0000000000000000", 26399 => "0000000000000000", 26400 => "0000000000000000", 26401 => "0000000000000000", 26402 => "0000000000000000", 26403 => "0000000000000000", 26404 => "0000000000000000", 26405 => "0000000000000000", 26406 => "0000000000000000", 26407 => "0000000000000000", 26408 => "0000000000000000", 26409 => "0000000000000000", 26410 => "0000000000000000", 26411 => "0000000000000000", 26412 => "0000000000000000", 26413 => "0000000000000000", 26414 => "0000000000000000", 26415 => "0000000000000000", 26416 => "0000000000000000", 26417 => "0000000000000000", 26418 => "0000000000000000", 26419 => "0000000000000000", 26420 => "0000000000000000", 26421 => "0000000000000000", 26422 => "0000000000000000", 26423 => "0000000000000000", 26424 => "0000000000000000", 26425 => "0000000000000000", 26426 => "0000000000000000", 26427 => "0000000000000000", 26428 => "0000000000000000", 26429 => "0000000000000000", 26430 => "0000000000000000", 26431 => "0000000000000000", 26432 => "0000000000000000", 26433 => "0000000000000000", 26434 => "0000000000000000", 26435 => "0000000000000000", 26436 => "0000000000000000", 26437 => "0000000000000000", 26438 => "0000000000000000", 26439 => "0000000000000000", 26440 => "0000000000000000", 26441 => "0000000000000000", 26442 => "0000000000000000", 26443 => "0000000000000000", 26444 => "0000000000000000", 26445 => "0000000000000000", 26446 => "0000000000000000", 26447 => "0000000000000000", 26448 => "0000000000000000", 26449 => "0000000000000000", 26450 => "0000000000000000", 26451 => "0000000000000000", 26452 => "0000000000000000", 26453 => "0000000000000000", 26454 => "0000000000000000", 26455 => "0000000000000000", 26456 => "0000000000000000", 26457 => "0000000000000000", 26458 => "0000000000000000", 26459 => "0000000000000000", 26460 => "0000000000000000", 26461 => "0000000000000000", 26462 => "0000000000000000", 26463 => "0000000000000000", 26464 => "0000000000000000", 26465 => "0000000000000000", 26466 => "0000000000000000", 26467 => "0000000000000000", 26468 => "0000000000000000", 26469 => "0000000000000000", 26470 => "0000000000000000", 26471 => "0000000000000000", 26472 => "0000000000000000", 26473 => "0000000000000000", 26474 => "0000000000000000", 26475 => "0000000000000000", 26476 => "0000000000000000", 26477 => "0000000000000000", 26478 => "0000000000000000", 26479 => "0000000000000000", 26480 => "0000000000000000", 26481 => "0000000000000000", 26482 => "0000000000000000", 26483 => "0000000000000000", 26484 => "0000000000000000", 26485 => "0000000000000000", 26486 => "0000000000000000", 26487 => "0000000000000000", 26488 => "0000000000000000", 26489 => "0000000000000000", 26490 => "0000000000000000", 26491 => "0000000000000000", 26492 => "0000000000000000", 26493 => "0000000000000000", 26494 => "0000000000000000", 26495 => "0000000000000000", 26496 => "0000000000000000", 26497 => "0000000000000000", 26498 => "0000000000000000", 26499 => "0000000000000000", 26500 => "0000000000000000", 26501 => "0000000000000000", 26502 => "0000000000000000", 26503 => "0000000000000000", 26504 => "0000000000000000", 26505 => "0000000000000000", 26506 => "0000000000000000", 26507 => "0000000000000000", 26508 => "0000000000000000", 26509 => "0000000000000000", 26510 => "0000000000000000", 26511 => "0000000000000000", 26512 => "0000000000000000", 26513 => "0000000000000000", 26514 => "0000000000000000", 26515 => "0000000000000000", 26516 => "0000000000000000", 26517 => "0000000000000000", 26518 => "0000000000000000", 26519 => "0000000000000000", 26520 => "0000000000000000", 26521 => "0000000000000000", 26522 => "0000000000000000", 26523 => "0000000000000000", 26524 => "0000000000000000", 26525 => "0000000000000000", 26526 => "0000000000000000", 26527 => "0000000000000000", 26528 => "0000000000000000", 26529 => "0000000000000000", 26530 => "0000000000000000", 26531 => "0000000000000000", 26532 => "0000000000000000", 26533 => "0000000000000000", 26534 => "0000000000000000", 26535 => "0000000000000000", 26536 => "0000000000000000", 26537 => "0000000000000000", 26538 => "0000000000000000", 26539 => "0000000000000000", 26540 => "0000000000000000", 26541 => "0000000000000000", 26542 => "0000000000000000", 26543 => "0000000000000000", 26544 => "0000000000000000", 26545 => "0000000000000000", 26546 => "0000000000000000", 26547 => "0000000000000000", 26548 => "0000000000000000", 26549 => "0000000000000000", 26550 => "0000000000000000", 26551 => "0000000000000000", 26552 => "0000000000000000", 26553 => "0000000000000000", 26554 => "0000000000000000", 26555 => "0000000000000000", 26556 => "0000000000000000", 26557 => "0000000000000000", 26558 => "0000000000000000", 26559 => "0000000000000000", 26560 => "0000000000000000", 26561 => "0000000000000000", 26562 => "0000000000000000", 26563 => "0000000000000000", 26564 => "0000000000000000", 26565 => "0000000000000000", 26566 => "0000000000000000", 26567 => "0000000000000000", 26568 => "0000000000000000", 26569 => "0000000000000000", 26570 => "0000000000000000", 26571 => "0000000000000000", 26572 => "0000000000000000", 26573 => "0000000000000000", 26574 => "0000000000000000", 26575 => "0000000000000000", 26576 => "0000000000000000", 26577 => "0000000000000000", 26578 => "0000000000000000", 26579 => "0000000000000000", 26580 => "0000000000000000", 26581 => "0000000000000000", 26582 => "0000000000000000", 26583 => "0000000000000000", 26584 => "0000000000000000", 26585 => "0000000000000000", 26586 => "0000000000000000", 26587 => "0000000000000000", 26588 => "0000000000000000", 26589 => "0000000000000000", 26590 => "0000000000000000", 26591 => "0000000000000000", 26592 => "0000000000000000", 26593 => "0000000000000000", 26594 => "0000000000000000", 26595 => "0000000000000000", 26596 => "0000000000000000", 26597 => "0000000000000000", 26598 => "0000000000000000", 26599 => "0000000000000000", 26600 => "0000000000000000", 26601 => "0000000000000000", 26602 => "0000000000000000", 26603 => "0000000000000000", 26604 => "0000000000000000", 26605 => "0000000000000000", 26606 => "0000000000000000", 26607 => "0000000000000000", 26608 => "0000000000000000", 26609 => "0000000000000000", 26610 => "0000000000000000", 26611 => "0000000000000000", 26612 => "0000000000000000", 26613 => "0000000000000000", 26614 => "0000000000000000", 26615 => "0000000000000000", 26616 => "0000000000000000", 26617 => "0000000000000000", 26618 => "0000000000000000", 26619 => "0000000000000000", 26620 => "0000000000000000", 26621 => "0000000000000000", 26622 => "0000000000000000", 26623 => "0000000000000000", 26624 => "0000000000000000", 26625 => "0000000000000000", 26626 => "0000000000000000", 26627 => "0000000000000000", 26628 => "0000000000000000", 26629 => "0000000000000000", 26630 => "0000000000000000", 26631 => "0000000000000000", 26632 => "0000000000000000", 26633 => "0000000000000000", 26634 => "0000000000000000", 26635 => "0000000000000000", 26636 => "0000000000000000", 26637 => "0000000000000000", 26638 => "0000000000000000", 26639 => "0000000000000000", 26640 => "0000000000000000", 26641 => "0000000000000000", 26642 => "0000000000000000", 26643 => "0000000000000000", 26644 => "0000000000000000", 26645 => "0000000000000000", 26646 => "0000000000000000", 26647 => "0000000000000000", 26648 => "0000000000000000", 26649 => "0000000000000000", 26650 => "0000000000000000", 26651 => "0000000000000000", 26652 => "0000000000000000", 26653 => "0000000000000000", 26654 => "0000000000000000", 26655 => "0000000000000000", 26656 => "0000000000000000", 26657 => "0000000000000000", 26658 => "0000000000000000", 26659 => "0000000000000000", 26660 => "0000000000000000", 26661 => "0000000000000000", 26662 => "0000000000000000", 26663 => "0000000000000000", 26664 => "0000000000000000", 26665 => "0000000000000000", 26666 => "0000000000000000", 26667 => "0000000000000000", 26668 => "0000000000000000", 26669 => "0000000000000000", 26670 => "0000000000000000", 26671 => "0000000000000000", 26672 => "0000000000000000", 26673 => "0000000000000000", 26674 => "0000000000000000", 26675 => "0000000000000000", 26676 => "0000000000000000", 26677 => "0000000000000000", 26678 => "0000000000000000", 26679 => "0000000000000000", 26680 => "0000000000000000", 26681 => "0000000000000000", 26682 => "0000000000000000", 26683 => "0000000000000000", 26684 => "0000000000000000", 26685 => "0000000000000000", 26686 => "0000000000000000", 26687 => "0000000000000000", 26688 => "0000000000000000", 26689 => "0000000000000000", 26690 => "0000000000000000", 26691 => "0000000000000000", 26692 => "0000000000000000", 26693 => "0000000000000000", 26694 => "0000000000000000", 26695 => "0000000000000000", 26696 => "0000000000000000", 26697 => "0000000000000000", 26698 => "0000000000000000", 26699 => "0000000000000000", 26700 => "0000000000000000", 26701 => "0000000000000000", 26702 => "0000000000000000", 26703 => "0000000000000000", 26704 => "0000000000000000", 26705 => "0000000000000000", 26706 => "0000000000000000", 26707 => "0000000000000000", 26708 => "0000000000000000", 26709 => "0000000000000000", 26710 => "0000000000000000", 26711 => "0000000000000000", 26712 => "0000000000000000", 26713 => "0000000000000000", 26714 => "0000000000000000", 26715 => "0000000000000000", 26716 => "0000000000000000", 26717 => "0000000000000000", 26718 => "0000000000000000", 26719 => "0000000000000000", 26720 => "0000000000000000", 26721 => "0000000000000000", 26722 => "0000000000000000", 26723 => "0000000000000000", 26724 => "0000000000000000", 26725 => "0000000000000000", 26726 => "0000000000000000", 26727 => "0000000000000000", 26728 => "0000000000000000", 26729 => "0000000000000000", 26730 => "0000000000000000", 26731 => "0000000000000000", 26732 => "0000000000000000", 26733 => "0000000000000000", 26734 => "0000000000000000", 26735 => "0000000000000000", 26736 => "0000000000000000", 26737 => "0000000000000000", 26738 => "0000000000000000", 26739 => "0000000000000000", 26740 => "0000000000000000", 26741 => "0000000000000000", 26742 => "0000000000000000", 26743 => "0000000000000000", 26744 => "0000000000000000", 26745 => "0000000000000000", 26746 => "0000000000000000", 26747 => "0000000000000000", 26748 => "0000000000000000", 26749 => "0000000000000000", 26750 => "0000000000000000", 26751 => "0000000000000000", 26752 => "0000000000000000", 26753 => "0000000000000000", 26754 => "0000000000000000", 26755 => "0000000000000000", 26756 => "0000000000000000", 26757 => "0000000000000000", 26758 => "0000000000000000", 26759 => "0000000000000000", 26760 => "0000000000000000", 26761 => "0000000000000000", 26762 => "0000000000000000", 26763 => "0000000000000000", 26764 => "0000000000000000", 26765 => "0000000000000000", 26766 => "0000000000000000", 26767 => "0000000000000000", 26768 => "0000000000000000", 26769 => "0000000000000000", 26770 => "0000000000000000", 26771 => "0000000000000000", 26772 => "0000000000000000", 26773 => "0000000000000000", 26774 => "0000000000000000", 26775 => "0000000000000000", 26776 => "0000000000000000", 26777 => "0000000000000000", 26778 => "0000000000000000", 26779 => "0000000000000000", 26780 => "0000000000000000", 26781 => "0000000000000000", 26782 => "0000000000000000", 26783 => "0000000000000000", 26784 => "0000000000000000", 26785 => "0000000000000000", 26786 => "0000000000000000", 26787 => "0000000000000000", 26788 => "0000000000000000", 26789 => "0000000000000000", 26790 => "0000000000000000", 26791 => "0000000000000000", 26792 => "0000000000000000", 26793 => "0000000000000000", 26794 => "0000000000000000", 26795 => "0000000000000000", 26796 => "0000000000000000", 26797 => "0000000000000000", 26798 => "0000000000000000", 26799 => "0000000000000000", 26800 => "0000000000000000", 26801 => "0000000000000000", 26802 => "0000000000000000", 26803 => "0000000000000000", 26804 => "0000000000000000", 26805 => "0000000000000000", 26806 => "0000000000000000", 26807 => "0000000000000000", 26808 => "0000000000000000", 26809 => "0000000000000000", 26810 => "0000000000000000", 26811 => "0000000000000000", 26812 => "0000000000000000", 26813 => "0000000000000000", 26814 => "0000000000000000", 26815 => "0000000000000000", 26816 => "0000000000000000", 26817 => "0000000000000000", 26818 => "0000000000000000", 26819 => "0000000000000000", 26820 => "0000000000000000", 26821 => "0000000000000000", 26822 => "0000000000000000", 26823 => "0000000000000000", 26824 => "0000000000000000", 26825 => "0000000000000000", 26826 => "0000000000000000", 26827 => "0000000000000000", 26828 => "0000000000000000", 26829 => "0000000000000000", 26830 => "0000000000000000", 26831 => "0000000000000000", 26832 => "0000000000000000", 26833 => "0000000000000000", 26834 => "0000000000000000", 26835 => "0000000000000000", 26836 => "0000000000000000", 26837 => "0000000000000000", 26838 => "0000000000000000", 26839 => "0000000000000000", 26840 => "0000000000000000", 26841 => "0000000000000000", 26842 => "0000000000000000", 26843 => "0000000000000000", 26844 => "0000000000000000", 26845 => "0000000000000000", 26846 => "0000000000000000", 26847 => "0000000000000000", 26848 => "0000000000000000", 26849 => "0000000000000000", 26850 => "0000000000000000", 26851 => "0000000000000000", 26852 => "0000000000000000", 26853 => "0000000000000000", 26854 => "0000000000000000", 26855 => "0000000000000000", 26856 => "0000000000000000", 26857 => "0000000000000000", 26858 => "0000000000000000", 26859 => "0000000000000000", 26860 => "0000000000000000", 26861 => "0000000000000000", 26862 => "0000000000000000", 26863 => "0000000000000000", 26864 => "0000000000000000", 26865 => "0000000000000000", 26866 => "0000000000000000", 26867 => "0000000000000000", 26868 => "0000000000000000", 26869 => "0000000000000000", 26870 => "0000000000000000", 26871 => "0000000000000000", 26872 => "0000000000000000", 26873 => "0000000000000000", 26874 => "0000000000000000", 26875 => "0000000000000000", 26876 => "0000000000000000", 26877 => "0000000000000000", 26878 => "0000000000000000", 26879 => "0000000000000000", 26880 => "0000000000000000", 26881 => "0000000000000000", 26882 => "0000000000000000", 26883 => "0000000000000000", 26884 => "0000000000000000", 26885 => "0000000000000000", 26886 => "0000000000000000", 26887 => "0000000000000000", 26888 => "0000000000000000", 26889 => "0000000000000000", 26890 => "0000000000000000", 26891 => "0000000000000000", 26892 => "0000000000000000", 26893 => "0000000000000000", 26894 => "0000000000000000", 26895 => "0000000000000000", 26896 => "0000000000000000", 26897 => "0000000000000000", 26898 => "0000000000000000", 26899 => "0000000000000000", 26900 => "0000000000000000", 26901 => "0000000000000000", 26902 => "0000000000000000", 26903 => "0000000000000000", 26904 => "0000000000000000", 26905 => "0000000000000000", 26906 => "0000000000000000", 26907 => "0000000000000000", 26908 => "0000000000000000", 26909 => "0000000000000000", 26910 => "0000000000000000", 26911 => "0000000000000000", 26912 => "0000000000000000", 26913 => "0000000000000000", 26914 => "0000000000000000", 26915 => "0000000000000000", 26916 => "0000000000000000", 26917 => "0000000000000000", 26918 => "0000000000000000", 26919 => "0000000000000000", 26920 => "0000000000000000", 26921 => "0000000000000000", 26922 => "0000000000000000", 26923 => "0000000000000000", 26924 => "0000000000000000", 26925 => "0000000000000000", 26926 => "0000000000000000", 26927 => "0000000000000000", 26928 => "0000000000000000", 26929 => "0000000000000000", 26930 => "0000000000000000", 26931 => "0000000000000000", 26932 => "0000000000000000", 26933 => "0000000000000000", 26934 => "0000000000000000", 26935 => "0000000000000000", 26936 => "0000000000000000", 26937 => "0000000000000000", 26938 => "0000000000000000", 26939 => "0000000000000000", 26940 => "0000000000000000", 26941 => "0000000000000000", 26942 => "0000000000000000", 26943 => "0000000000000000", 26944 => "0000000000000000", 26945 => "0000000000000000", 26946 => "0000000000000000", 26947 => "0000000000000000", 26948 => "0000000000000000", 26949 => "0000000000000000", 26950 => "0000000000000000", 26951 => "0000000000000000", 26952 => "0000000000000000", 26953 => "0000000000000000", 26954 => "0000000000000000", 26955 => "0000000000000000", 26956 => "0000000000000000", 26957 => "0000000000000000", 26958 => "0000000000000000", 26959 => "0000000000000000", 26960 => "0000000000000000", 26961 => "0000000000000000", 26962 => "0000000000000000", 26963 => "0000000000000000", 26964 => "0000000000000000", 26965 => "0000000000000000", 26966 => "0000000000000000", 26967 => "0000000000000000", 26968 => "0000000000000000", 26969 => "0000000000000000", 26970 => "0000000000000000", 26971 => "0000000000000000", 26972 => "0000000000000000", 26973 => "0000000000000000", 26974 => "0000000000000000", 26975 => "0000000000000000", 26976 => "0000000000000000", 26977 => "0000000000000000", 26978 => "0000000000000000", 26979 => "0000000000000000", 26980 => "0000000000000000", 26981 => "0000000000000000", 26982 => "0000000000000000", 26983 => "0000000000000000", 26984 => "0000000000000000", 26985 => "0000000000000000", 26986 => "0000000000000000", 26987 => "0000000000000000", 26988 => "0000000000000000", 26989 => "0000000000000000", 26990 => "0000000000000000", 26991 => "0000000000000000", 26992 => "0000000000000000", 26993 => "0000000000000000", 26994 => "0000000000000000", 26995 => "0000000000000000", 26996 => "0000000000000000", 26997 => "0000000000000000", 26998 => "0000000000000000", 26999 => "0000000000000000", 27000 => "0000000000000000", 27001 => "0000000000000000", 27002 => "0000000000000000", 27003 => "0000000000000000", 27004 => "0000000000000000", 27005 => "0000000000000000", 27006 => "0000000000000000", 27007 => "0000000000000000", 27008 => "0000000000000000", 27009 => "0000000000000000", 27010 => "0000000000000000", 27011 => "0000000000000000", 27012 => "0000000000000000", 27013 => "0000000000000000", 27014 => "0000000000000000", 27015 => "0000000000000000", 27016 => "0000000000000000", 27017 => "0000000000000000", 27018 => "0000000000000000", 27019 => "0000000000000000", 27020 => "0000000000000000", 27021 => "0000000000000000", 27022 => "0000000000000000", 27023 => "0000000000000000", 27024 => "0000000000000000", 27025 => "0000000000000000", 27026 => "0000000000000000", 27027 => "0000000000000000", 27028 => "0000000000000000", 27029 => "0000000000000000", 27030 => "0000000000000000", 27031 => "0000000000000000", 27032 => "0000000000000000", 27033 => "0000000000000000", 27034 => "0000000000000000", 27035 => "0000000000000000", 27036 => "0000000000000000", 27037 => "0000000000000000", 27038 => "0000000000000000", 27039 => "0000000000000000", 27040 => "0000000000000000", 27041 => "0000000000000000", 27042 => "0000000000000000", 27043 => "0000000000000000", 27044 => "0000000000000000", 27045 => "0000000000000000", 27046 => "0000000000000000", 27047 => "0000000000000000", 27048 => "0000000000000000", 27049 => "0000000000000000", 27050 => "0000000000000000", 27051 => "0000000000000000", 27052 => "0000000000000000", 27053 => "0000000000000000", 27054 => "0000000000000000", 27055 => "0000000000000000", 27056 => "0000000000000000", 27057 => "0000000000000000", 27058 => "0000000000000000", 27059 => "0000000000000000", 27060 => "0000000000000000", 27061 => "0000000000000000", 27062 => "0000000000000000", 27063 => "0000000000000000", 27064 => "0000000000000000", 27065 => "0000000000000000", 27066 => "0000000000000000", 27067 => "0000000000000000", 27068 => "0000000000000000", 27069 => "0000000000000000", 27070 => "0000000000000000", 27071 => "0000000000000000", 27072 => "0000000000000000", 27073 => "0000000000000000", 27074 => "0000000000000000", 27075 => "0000000000000000", 27076 => "0000000000000000", 27077 => "0000000000000000", 27078 => "0000000000000000", 27079 => "0000000000000000", 27080 => "0000000000000000", 27081 => "0000000000000000", 27082 => "0000000000000000", 27083 => "0000000000000000", 27084 => "0000000000000000", 27085 => "0000000000000000", 27086 => "0000000000000000", 27087 => "0000000000000000", 27088 => "0000000000000000", 27089 => "0000000000000000", 27090 => "0000000000000000", 27091 => "0000000000000000", 27092 => "0000000000000000", 27093 => "0000000000000000", 27094 => "0000000000000000", 27095 => "0000000000000000", 27096 => "0000000000000000", 27097 => "0000000000000000", 27098 => "0000000000000000", 27099 => "0000000000000000", 27100 => "0000000000000000", 27101 => "0000000000000000", 27102 => "0000000000000000", 27103 => "0000000000000000", 27104 => "0000000000000000", 27105 => "0000000000000000", 27106 => "0000000000000000", 27107 => "0000000000000000", 27108 => "0000000000000000", 27109 => "0000000000000000", 27110 => "0000000000000000", 27111 => "0000000000000000", 27112 => "0000000000000000", 27113 => "0000000000000000", 27114 => "0000000000000000", 27115 => "0000000000000000", 27116 => "0000000000000000", 27117 => "0000000000000000", 27118 => "0000000000000000", 27119 => "0000000000000000", 27120 => "0000000000000000", 27121 => "0000000000000000", 27122 => "0000000000000000", 27123 => "0000000000000000", 27124 => "0000000000000000", 27125 => "0000000000000000", 27126 => "0000000000000000", 27127 => "0000000000000000", 27128 => "0000000000000000", 27129 => "0000000000000000", 27130 => "0000000000000000", 27131 => "0000000000000000", 27132 => "0000000000000000", 27133 => "0000000000000000", 27134 => "0000000000000000", 27135 => "0000000000000000", 27136 => "0000000000000000", 27137 => "0000000000000000", 27138 => "0000000000000000", 27139 => "0000000000000000", 27140 => "0000000000000000", 27141 => "0000000000000000", 27142 => "0000000000000000", 27143 => "0000000000000000", 27144 => "0000000000000000", 27145 => "0000000000000000", 27146 => "0000000000000000", 27147 => "0000000000000000", 27148 => "0000000000000000", 27149 => "0000000000000000", 27150 => "0000000000000000", 27151 => "0000000000000000", 27152 => "0000000000000000", 27153 => "0000000000000000", 27154 => "0000000000000000", 27155 => "0000000000000000", 27156 => "0000000000000000", 27157 => "0000000000000000", 27158 => "0000000000000000", 27159 => "0000000000000000", 27160 => "0000000000000000", 27161 => "0000000000000000", 27162 => "0000000000000000", 27163 => "0000000000000000", 27164 => "0000000000000000", 27165 => "0000000000000000", 27166 => "0000000000000000", 27167 => "0000000000000000", 27168 => "0000000000000000", 27169 => "0000000000000000", 27170 => "0000000000000000", 27171 => "0000000000000000", 27172 => "0000000000000000", 27173 => "0000000000000000", 27174 => "0000000000000000", 27175 => "0000000000000000", 27176 => "0000000000000000", 27177 => "0000000000000000", 27178 => "0000000000000000", 27179 => "0000000000000000", 27180 => "0000000000000000", 27181 => "0000000000000000", 27182 => "0000000000000000", 27183 => "0000000000000000", 27184 => "0000000000000000", 27185 => "0000000000000000", 27186 => "0000000000000000", 27187 => "0000000000000000", 27188 => "0000000000000000", 27189 => "0000000000000000", 27190 => "0000000000000000", 27191 => "0000000000000000", 27192 => "0000000000000000", 27193 => "0000000000000000", 27194 => "0000000000000000", 27195 => "0000000000000000", 27196 => "0000000000000000", 27197 => "0000000000000000", 27198 => "0000000000000000", 27199 => "0000000000000000", 27200 => "0000000000000000", 27201 => "0000000000000000", 27202 => "0000000000000000", 27203 => "0000000000000000", 27204 => "0000000000000000", 27205 => "0000000000000000", 27206 => "0000000000000000", 27207 => "0000000000000000", 27208 => "0000000000000000", 27209 => "0000000000000000", 27210 => "0000000000000000", 27211 => "0000000000000000", 27212 => "0000000000000000", 27213 => "0000000000000000", 27214 => "0000000000000000", 27215 => "0000000000000000", 27216 => "0000000000000000", 27217 => "0000000000000000", 27218 => "0000000000000000", 27219 => "0000000000000000", 27220 => "0000000000000000", 27221 => "0000000000000000", 27222 => "0000000000000000", 27223 => "0000000000000000", 27224 => "0000000000000000", 27225 => "0000000000000000", 27226 => "0000000000000000", 27227 => "0000000000000000", 27228 => "0000000000000000", 27229 => "0000000000000000", 27230 => "0000000000000000", 27231 => "0000000000000000", 27232 => "0000000000000000", 27233 => "0000000000000000", 27234 => "0000000000000000", 27235 => "0000000000000000", 27236 => "0000000000000000", 27237 => "0000000000000000", 27238 => "0000000000000000", 27239 => "0000000000000000", 27240 => "0000000000000000", 27241 => "0000000000000000", 27242 => "0000000000000000", 27243 => "0000000000000000", 27244 => "0000000000000000", 27245 => "0000000000000000", 27246 => "0000000000000000", 27247 => "0000000000000000", 27248 => "0000000000000000", 27249 => "0000000000000000", 27250 => "0000000000000000", 27251 => "0000000000000000", 27252 => "0000000000000000", 27253 => "0000000000000000", 27254 => "0000000000000000", 27255 => "0000000000000000", 27256 => "0000000000000000", 27257 => "0000000000000000", 27258 => "0000000000000000", 27259 => "0000000000000000", 27260 => "0000000000000000", 27261 => "0000000000000000", 27262 => "0000000000000000", 27263 => "0000000000000000", 27264 => "0000000000000000", 27265 => "0000000000000000", 27266 => "0000000000000000", 27267 => "0000000000000000", 27268 => "0000000000000000", 27269 => "0000000000000000", 27270 => "0000000000000000", 27271 => "0000000000000000", 27272 => "0000000000000000", 27273 => "0000000000000000", 27274 => "0000000000000000", 27275 => "0000000000000000", 27276 => "0000000000000000", 27277 => "0000000000000000", 27278 => "0000000000000000", 27279 => "0000000000000000", 27280 => "0000000000000000", 27281 => "0000000000000000", 27282 => "0000000000000000", 27283 => "0000000000000000", 27284 => "0000000000000000", 27285 => "0000000000000000", 27286 => "0000000000000000", 27287 => "0000000000000000", 27288 => "0000000000000000", 27289 => "0000000000000000", 27290 => "0000000000000000", 27291 => "0000000000000000", 27292 => "0000000000000000", 27293 => "0000000000000000", 27294 => "0000000000000000", 27295 => "0000000000000000", 27296 => "0000000000000000", 27297 => "0000000000000000", 27298 => "0000000000000000", 27299 => "0000000000000000", 27300 => "0000000000000000", 27301 => "0000000000000000", 27302 => "0000000000000000", 27303 => "0000000000000000", 27304 => "0000000000000000", 27305 => "0000000000000000", 27306 => "0000000000000000", 27307 => "0000000000000000", 27308 => "0000000000000000", 27309 => "0000000000000000", 27310 => "0000000000000000", 27311 => "0000000000000000", 27312 => "0000000000000000", 27313 => "0000000000000000", 27314 => "0000000000000000", 27315 => "0000000000000000", 27316 => "0000000000000000", 27317 => "0000000000000000", 27318 => "0000000000000000", 27319 => "0000000000000000", 27320 => "0000000000000000", 27321 => "0000000000000000", 27322 => "0000000000000000", 27323 => "0000000000000000", 27324 => "0000000000000000", 27325 => "0000000000000000", 27326 => "0000000000000000", 27327 => "0000000000000000", 27328 => "0000000000000000", 27329 => "0000000000000000", 27330 => "0000000000000000", 27331 => "0000000000000000", 27332 => "0000000000000000", 27333 => "0000000000000000", 27334 => "0000000000000000", 27335 => "0000000000000000", 27336 => "0000000000000000", 27337 => "0000000000000000", 27338 => "0000000000000000", 27339 => "0000000000000000", 27340 => "0000000000000000", 27341 => "0000000000000000", 27342 => "0000000000000000", 27343 => "0000000000000000", 27344 => "0000000000000000", 27345 => "0000000000000000", 27346 => "0000000000000000", 27347 => "0000000000000000", 27348 => "0000000000000000", 27349 => "0000000000000000", 27350 => "0000000000000000", 27351 => "0000000000000000", 27352 => "0000000000000000", 27353 => "0000000000000000", 27354 => "0000000000000000", 27355 => "0000000000000000", 27356 => "0000000000000000", 27357 => "0000000000000000", 27358 => "0000000000000000", 27359 => "0000000000000000", 27360 => "0000000000000000", 27361 => "0000000000000000", 27362 => "0000000000000000", 27363 => "0000000000000000", 27364 => "0000000000000000", 27365 => "0000000000000000", 27366 => "0000000000000000", 27367 => "0000000000000000", 27368 => "0000000000000000", 27369 => "0000000000000000", 27370 => "0000000000000000", 27371 => "0000000000000000", 27372 => "0000000000000000", 27373 => "0000000000000000", 27374 => "0000000000000000", 27375 => "0000000000000000", 27376 => "0000000000000000", 27377 => "0000000000000000", 27378 => "0000000000000000", 27379 => "0000000000000000", 27380 => "0000000000000000", 27381 => "0000000000000000", 27382 => "0000000000000000", 27383 => "0000000000000000", 27384 => "0000000000000000", 27385 => "0000000000000000", 27386 => "0000000000000000", 27387 => "0000000000000000", 27388 => "0000000000000000", 27389 => "0000000000000000", 27390 => "0000000000000000", 27391 => "0000000000000000", 27392 => "0000000000000000", 27393 => "0000000000000000", 27394 => "0000000000000000", 27395 => "0000000000000000", 27396 => "0000000000000000", 27397 => "0000000000000000", 27398 => "0000000000000000", 27399 => "0000000000000000", 27400 => "0000000000000000", 27401 => "0000000000000000", 27402 => "0000000000000000", 27403 => "0000000000000000", 27404 => "0000000000000000", 27405 => "0000000000000000", 27406 => "0000000000000000", 27407 => "0000000000000000", 27408 => "0000000000000000", 27409 => "0000000000000000", 27410 => "0000000000000000", 27411 => "0000000000000000", 27412 => "0000000000000000", 27413 => "0000000000000000", 27414 => "0000000000000000", 27415 => "0000000000000000", 27416 => "0000000000000000", 27417 => "0000000000000000", 27418 => "0000000000000000", 27419 => "0000000000000000", 27420 => "0000000000000000", 27421 => "0000000000000000", 27422 => "0000000000000000", 27423 => "0000000000000000", 27424 => "0000000000000000", 27425 => "0000000000000000", 27426 => "0000000000000000", 27427 => "0000000000000000", 27428 => "0000000000000000", 27429 => "0000000000000000", 27430 => "0000000000000000", 27431 => "0000000000000000", 27432 => "0000000000000000", 27433 => "0000000000000000", 27434 => "0000000000000000", 27435 => "0000000000000000", 27436 => "0000000000000000", 27437 => "0000000000000000", 27438 => "0000000000000000", 27439 => "0000000000000000", 27440 => "0000000000000000", 27441 => "0000000000000000", 27442 => "0000000000000000", 27443 => "0000000000000000", 27444 => "0000000000000000", 27445 => "0000000000000000", 27446 => "0000000000000000", 27447 => "0000000000000000", 27448 => "0000000000000000", 27449 => "0000000000000000", 27450 => "0000000000000000", 27451 => "0000000000000000", 27452 => "0000000000000000", 27453 => "0000000000000000", 27454 => "0000000000000000", 27455 => "0000000000000000", 27456 => "0000000000000000", 27457 => "0000000000000000", 27458 => "0000000000000000", 27459 => "0000000000000000", 27460 => "0000000000000000", 27461 => "0000000000000000", 27462 => "0000000000000000", 27463 => "0000000000000000", 27464 => "0000000000000000", 27465 => "0000000000000000", 27466 => "0000000000000000", 27467 => "0000000000000000", 27468 => "0000000000000000", 27469 => "0000000000000000", 27470 => "0000000000000000", 27471 => "0000000000000000", 27472 => "0000000000000000", 27473 => "0000000000000000", 27474 => "0000000000000000", 27475 => "0000000000000000", 27476 => "0000000000000000", 27477 => "0000000000000000", 27478 => "0000000000000000", 27479 => "0000000000000000", 27480 => "0000000000000000", 27481 => "0000000000000000", 27482 => "0000000000000000", 27483 => "0000000000000000", 27484 => "0000000000000000", 27485 => "0000000000000000", 27486 => "0000000000000000", 27487 => "0000000000000000", 27488 => "0000000000000000", 27489 => "0000000000000000", 27490 => "0000000000000000", 27491 => "0000000000000000", 27492 => "0000000000000000", 27493 => "0000000000000000", 27494 => "0000000000000000", 27495 => "0000000000000000", 27496 => "0000000000000000", 27497 => "0000000000000000", 27498 => "0000000000000000", 27499 => "0000000000000000", 27500 => "0000000000000000", 27501 => "0000000000000000", 27502 => "0000000000000000", 27503 => "0000000000000000", 27504 => "0000000000000000", 27505 => "0000000000000000", 27506 => "0000000000000000", 27507 => "0000000000000000", 27508 => "0000000000000000", 27509 => "0000000000000000", 27510 => "0000000000000000", 27511 => "0000000000000000", 27512 => "0000000000000000", 27513 => "0000000000000000", 27514 => "0000000000000000", 27515 => "0000000000000000", 27516 => "0000000000000000", 27517 => "0000000000000000", 27518 => "0000000000000000", 27519 => "0000000000000000", 27520 => "0000000000000000", 27521 => "0000000000000000", 27522 => "0000000000000000", 27523 => "0000000000000000", 27524 => "0000000000000000", 27525 => "0000000000000000", 27526 => "0000000000000000", 27527 => "0000000000000000", 27528 => "0000000000000000", 27529 => "0000000000000000", 27530 => "0000000000000000", 27531 => "0000000000000000", 27532 => "0000000000000000", 27533 => "0000000000000000", 27534 => "0000000000000000", 27535 => "0000000000000000", 27536 => "0000000000000000", 27537 => "0000000000000000", 27538 => "0000000000000000", 27539 => "0000000000000000", 27540 => "0000000000000000", 27541 => "0000000000000000", 27542 => "0000000000000000", 27543 => "0000000000000000", 27544 => "0000000000000000", 27545 => "0000000000000000", 27546 => "0000000000000000", 27547 => "0000000000000000", 27548 => "0000000000000000", 27549 => "0000000000000000", 27550 => "0000000000000000", 27551 => "0000000000000000", 27552 => "0000000000000000", 27553 => "0000000000000000", 27554 => "0000000000000000", 27555 => "0000000000000000", 27556 => "0000000000000000", 27557 => "0000000000000000", 27558 => "0000000000000000", 27559 => "0000000000000000", 27560 => "0000000000000000", 27561 => "0000000000000000", 27562 => "0000000000000000", 27563 => "0000000000000000", 27564 => "0000000000000000", 27565 => "0000000000000000", 27566 => "0000000000000000", 27567 => "0000000000000000", 27568 => "0000000000000000", 27569 => "0000000000000000", 27570 => "0000000000000000", 27571 => "0000000000000000", 27572 => "0000000000000000", 27573 => "0000000000000000", 27574 => "0000000000000000", 27575 => "0000000000000000", 27576 => "0000000000000000", 27577 => "0000000000000000", 27578 => "0000000000000000", 27579 => "0000000000000000", 27580 => "0000000000000000", 27581 => "0000000000000000", 27582 => "0000000000000000", 27583 => "0000000000000000", 27584 => "0000000000000000", 27585 => "0000000000000000", 27586 => "0000000000000000", 27587 => "0000000000000000", 27588 => "0000000000000000", 27589 => "0000000000000000", 27590 => "0000000000000000", 27591 => "0000000000000000", 27592 => "0000000000000000", 27593 => "0000000000000000", 27594 => "0000000000000000", 27595 => "0000000000000000", 27596 => "0000000000000000", 27597 => "0000000000000000", 27598 => "0000000000000000", 27599 => "0000000000000000", 27600 => "0000000000000000", 27601 => "0000000000000000", 27602 => "0000000000000000", 27603 => "0000000000000000", 27604 => "0000000000000000", 27605 => "0000000000000000", 27606 => "0000000000000000", 27607 => "0000000000000000", 27608 => "0000000000000000", 27609 => "0000000000000000", 27610 => "0000000000000000", 27611 => "0000000000000000", 27612 => "0000000000000000", 27613 => "0000000000000000", 27614 => "0000000000000000", 27615 => "0000000000000000", 27616 => "0000000000000000", 27617 => "0000000000000000", 27618 => "0000000000000000", 27619 => "0000000000000000", 27620 => "0000000000000000", 27621 => "0000000000000000", 27622 => "0000000000000000", 27623 => "0000000000000000", 27624 => "0000000000000000", 27625 => "0000000000000000", 27626 => "0000000000000000", 27627 => "0000000000000000", 27628 => "0000000000000000", 27629 => "0000000000000000", 27630 => "0000000000000000", 27631 => "0000000000000000", 27632 => "0000000000000000", 27633 => "0000000000000000", 27634 => "0000000000000000", 27635 => "0000000000000000", 27636 => "0000000000000000", 27637 => "0000000000000000", 27638 => "0000000000000000", 27639 => "0000000000000000", 27640 => "0000000000000000", 27641 => "0000000000000000", 27642 => "0000000000000000", 27643 => "0000000000000000", 27644 => "0000000000000000", 27645 => "0000000000000000", 27646 => "0000000000000000", 27647 => "0000000000000000", 27648 => "0000000000000000", 27649 => "0000000000000000", 27650 => "0000000000000000", 27651 => "0000000000000000", 27652 => "0000000000000000", 27653 => "0000000000000000", 27654 => "0000000000000000", 27655 => "0000000000000000", 27656 => "0000000000000000", 27657 => "0000000000000000", 27658 => "0000000000000000", 27659 => "0000000000000000", 27660 => "0000000000000000", 27661 => "0000000000000000", 27662 => "0000000000000000", 27663 => "0000000000000000", 27664 => "0000000000000000", 27665 => "0000000000000000", 27666 => "0000000000000000", 27667 => "0000000000000000", 27668 => "0000000000000000", 27669 => "0000000000000000", 27670 => "0000000000000000", 27671 => "0000000000000000", 27672 => "0000000000000000", 27673 => "0000000000000000", 27674 => "0000000000000000", 27675 => "0000000000000000", 27676 => "0000000000000000", 27677 => "0000000000000000", 27678 => "0000000000000000", 27679 => "0000000000000000", 27680 => "0000000000000000", 27681 => "0000000000000000", 27682 => "0000000000000000", 27683 => "0000000000000000", 27684 => "0000000000000000", 27685 => "0000000000000000", 27686 => "0000000000000000", 27687 => "0000000000000000", 27688 => "0000000000000000", 27689 => "0000000000000000", 27690 => "0000000000000000", 27691 => "0000000000000000", 27692 => "0000000000000000", 27693 => "0000000000000000", 27694 => "0000000000000000", 27695 => "0000000000000000", 27696 => "0000000000000000", 27697 => "0000000000000000", 27698 => "0000000000000000", 27699 => "0000000000000000", 27700 => "0000000000000000", 27701 => "0000000000000000", 27702 => "0000000000000000", 27703 => "0000000000000000", 27704 => "0000000000000000", 27705 => "0000000000000000", 27706 => "0000000000000000", 27707 => "0000000000000000", 27708 => "0000000000000000", 27709 => "0000000000000000", 27710 => "0000000000000000", 27711 => "0000000000000000", 27712 => "0000000000000000", 27713 => "0000000000000000", 27714 => "0000000000000000", 27715 => "0000000000000000", 27716 => "0000000000000000", 27717 => "0000000000000000", 27718 => "0000000000000000", 27719 => "0000000000000000", 27720 => "0000000000000000", 27721 => "0000000000000000", 27722 => "0000000000000000", 27723 => "0000000000000000", 27724 => "0000000000000000", 27725 => "0000000000000000", 27726 => "0000000000000000", 27727 => "0000000000000000", 27728 => "0000000000000000", 27729 => "0000000000000000", 27730 => "0000000000000000", 27731 => "0000000000000000", 27732 => "0000000000000000", 27733 => "0000000000000000", 27734 => "0000000000000000", 27735 => "0000000000000000", 27736 => "0000000000000000", 27737 => "0000000000000000", 27738 => "0000000000000000", 27739 => "0000000000000000", 27740 => "0000000000000000", 27741 => "0000000000000000", 27742 => "0000000000000000", 27743 => "0000000000000000", 27744 => "0000000000000000", 27745 => "0000000000000000", 27746 => "0000000000000000", 27747 => "0000000000000000", 27748 => "0000000000000000", 27749 => "0000000000000000", 27750 => "0000000000000000", 27751 => "0000000000000000", 27752 => "0000000000000000", 27753 => "0000000000000000", 27754 => "0000000000000000", 27755 => "0000000000000000", 27756 => "0000000000000000", 27757 => "0000000000000000", 27758 => "0000000000000000", 27759 => "0000000000000000", 27760 => "0000000000000000", 27761 => "0000000000000000", 27762 => "0000000000000000", 27763 => "0000000000000000", 27764 => "0000000000000000", 27765 => "0000000000000000", 27766 => "0000000000000000", 27767 => "0000000000000000", 27768 => "0000000000000000", 27769 => "0000000000000000", 27770 => "0000000000000000", 27771 => "0000000000000000", 27772 => "0000000000000000", 27773 => "0000000000000000", 27774 => "0000000000000000", 27775 => "0000000000000000", 27776 => "0000000000000000", 27777 => "0000000000000000", 27778 => "0000000000000000", 27779 => "0000000000000000", 27780 => "0000000000000000", 27781 => "0000000000000000", 27782 => "0000000000000000", 27783 => "0000000000000000", 27784 => "0000000000000000", 27785 => "0000000000000000", 27786 => "0000000000000000", 27787 => "0000000000000000", 27788 => "0000000000000000", 27789 => "0000000000000000", 27790 => "0000000000000000", 27791 => "0000000000000000", 27792 => "0000000000000000", 27793 => "0000000000000000", 27794 => "0000000000000000", 27795 => "0000000000000000", 27796 => "0000000000000000", 27797 => "0000000000000000", 27798 => "0000000000000000", 27799 => "0000000000000000", 27800 => "0000000000000000", 27801 => "0000000000000000", 27802 => "0000000000000000", 27803 => "0000000000000000", 27804 => "0000000000000000", 27805 => "0000000000000000", 27806 => "0000000000000000", 27807 => "0000000000000000", 27808 => "0000000000000000", 27809 => "0000000000000000", 27810 => "0000000000000000", 27811 => "0000000000000000", 27812 => "0000000000000000", 27813 => "0000000000000000", 27814 => "0000000000000000", 27815 => "0000000000000000", 27816 => "0000000000000000", 27817 => "0000000000000000", 27818 => "0000000000000000", 27819 => "0000000000000000", 27820 => "0000000000000000", 27821 => "0000000000000000", 27822 => "0000000000000000", 27823 => "0000000000000000", 27824 => "0000000000000000", 27825 => "0000000000000000", 27826 => "0000000000000000", 27827 => "0000000000000000", 27828 => "0000000000000000", 27829 => "0000000000000000", 27830 => "0000000000000000", 27831 => "0000000000000000", 27832 => "0000000000000000", 27833 => "0000000000000000", 27834 => "0000000000000000", 27835 => "0000000000000000", 27836 => "0000000000000000", 27837 => "0000000000000000", 27838 => "0000000000000000", 27839 => "0000000000000000", 27840 => "0000000000000000", 27841 => "0000000000000000", 27842 => "0000000000000000", 27843 => "0000000000000000", 27844 => "0000000000000000", 27845 => "0000000000000000", 27846 => "0000000000000000", 27847 => "0000000000000000", 27848 => "0000000000000000", 27849 => "0000000000000000", 27850 => "0000000000000000", 27851 => "0000000000000000", 27852 => "0000000000000000", 27853 => "0000000000000000", 27854 => "0000000000000000", 27855 => "0000000000000000", 27856 => "0000000000000000", 27857 => "0000000000000000", 27858 => "0000000000000000", 27859 => "0000000000000000", 27860 => "0000000000000000", 27861 => "0000000000000000", 27862 => "0000000000000000", 27863 => "0000000000000000", 27864 => "0000000000000000", 27865 => "0000000000000000", 27866 => "0000000000000000", 27867 => "0000000000000000", 27868 => "0000000000000000", 27869 => "0000000000000000", 27870 => "0000000000000000", 27871 => "0000000000000000", 27872 => "0000000000000000", 27873 => "0000000000000000", 27874 => "0000000000000000", 27875 => "0000000000000000", 27876 => "0000000000000000", 27877 => "0000000000000000", 27878 => "0000000000000000", 27879 => "0000000000000000", 27880 => "0000000000000000", 27881 => "0000000000000000", 27882 => "0000000000000000", 27883 => "0000000000000000", 27884 => "0000000000000000", 27885 => "0000000000000000", 27886 => "0000000000000000", 27887 => "0000000000000000", 27888 => "0000000000000000", 27889 => "0000000000000000", 27890 => "0000000000000000", 27891 => "0000000000000000", 27892 => "0000000000000000", 27893 => "0000000000000000", 27894 => "0000000000000000", 27895 => "0000000000000000", 27896 => "0000000000000000", 27897 => "0000000000000000", 27898 => "0000000000000000", 27899 => "0000000000000000", 27900 => "0000000000000000", 27901 => "0000000000000000", 27902 => "0000000000000000", 27903 => "0000000000000000", 27904 => "0000000000000000", 27905 => "0000000000000000", 27906 => "0000000000000000", 27907 => "0000000000000000", 27908 => "0000000000000000", 27909 => "0000000000000000", 27910 => "0000000000000000", 27911 => "0000000000000000", 27912 => "0000000000000000", 27913 => "0000000000000000", 27914 => "0000000000000000", 27915 => "0000000000000000", 27916 => "0000000000000000", 27917 => "0000000000000000", 27918 => "0000000000000000", 27919 => "0000000000000000", 27920 => "0000000000000000", 27921 => "0000000000000000", 27922 => "0000000000000000", 27923 => "0000000000000000", 27924 => "0000000000000000", 27925 => "0000000000000000", 27926 => "0000000000000000", 27927 => "0000000000000000", 27928 => "0000000000000000", 27929 => "0000000000000000", 27930 => "0000000000000000", 27931 => "0000000000000000", 27932 => "0000000000000000", 27933 => "0000000000000000", 27934 => "0000000000000000", 27935 => "0000000000000000", 27936 => "0000000000000000", 27937 => "0000000000000000", 27938 => "0000000000000000", 27939 => "0000000000000000", 27940 => "0000000000000000", 27941 => "0000000000000000", 27942 => "0000000000000000", 27943 => "0000000000000000", 27944 => "0000000000000000", 27945 => "0000000000000000", 27946 => "0000000000000000", 27947 => "0000000000000000", 27948 => "0000000000000000", 27949 => "0000000000000000", 27950 => "0000000000000000", 27951 => "0000000000000000", 27952 => "0000000000000000", 27953 => "0000000000000000", 27954 => "0000000000000000", 27955 => "0000000000000000", 27956 => "0000000000000000", 27957 => "0000000000000000", 27958 => "0000000000000000", 27959 => "0000000000000000", 27960 => "0000000000000000", 27961 => "0000000000000000", 27962 => "0000000000000000", 27963 => "0000000000000000", 27964 => "0000000000000000", 27965 => "0000000000000000", 27966 => "0000000000000000", 27967 => "0000000000000000", 27968 => "0000000000000000", 27969 => "0000000000000000", 27970 => "0000000000000000", 27971 => "0000000000000000", 27972 => "0000000000000000", 27973 => "0000000000000000", 27974 => "0000000000000000", 27975 => "0000000000000000", 27976 => "0000000000000000", 27977 => "0000000000000000", 27978 => "0000000000000000", 27979 => "0000000000000000", 27980 => "0000000000000000", 27981 => "0000000000000000", 27982 => "0000000000000000", 27983 => "0000000000000000", 27984 => "0000000000000000", 27985 => "0000000000000000", 27986 => "0000000000000000", 27987 => "0000000000000000", 27988 => "0000000000000000", 27989 => "0000000000000000", 27990 => "0000000000000000", 27991 => "0000000000000000", 27992 => "0000000000000000", 27993 => "0000000000000000", 27994 => "0000000000000000", 27995 => "0000000000000000", 27996 => "0000000000000000", 27997 => "0000000000000000", 27998 => "0000000000000000", 27999 => "0000000000000000", 28000 => "0000000000000000", 28001 => "0000000000000000", 28002 => "0000000000000000", 28003 => "0000000000000000", 28004 => "0000000000000000", 28005 => "0000000000000000", 28006 => "0000000000000000", 28007 => "0000000000000000", 28008 => "0000000000000000", 28009 => "0000000000000000", 28010 => "0000000000000000", 28011 => "0000000000000000", 28012 => "0000000000000000", 28013 => "0000000000000000", 28014 => "0000000000000000", 28015 => "0000000000000000", 28016 => "0000000000000000", 28017 => "0000000000000000", 28018 => "0000000000000000", 28019 => "0000000000000000", 28020 => "0000000000000000", 28021 => "0000000000000000", 28022 => "0000000000000000", 28023 => "0000000000000000", 28024 => "0000000000000000", 28025 => "0000000000000000", 28026 => "0000000000000000", 28027 => "0000000000000000", 28028 => "0000000000000000", 28029 => "0000000000000000", 28030 => "0000000000000000", 28031 => "0000000000000000", 28032 => "0000000000000000", 28033 => "0000000000000000", 28034 => "0000000000000000", 28035 => "0000000000000000", 28036 => "0000000000000000", 28037 => "0000000000000000", 28038 => "0000000000000000", 28039 => "0000000000000000", 28040 => "0000000000000000", 28041 => "0000000000000000", 28042 => "0000000000000000", 28043 => "0000000000000000", 28044 => "0000000000000000", 28045 => "0000000000000000", 28046 => "0000000000000000", 28047 => "0000000000000000", 28048 => "0000000000000000", 28049 => "0000000000000000", 28050 => "0000000000000000", 28051 => "0000000000000000", 28052 => "0000000000000000", 28053 => "0000000000000000", 28054 => "0000000000000000", 28055 => "0000000000000000", 28056 => "0000000000000000", 28057 => "0000000000000000", 28058 => "0000000000000000", 28059 => "0000000000000000", 28060 => "0000000000000000", 28061 => "0000000000000000", 28062 => "0000000000000000", 28063 => "0000000000000000", 28064 => "0000000000000000", 28065 => "0000000000000000", 28066 => "0000000000000000", 28067 => "0000000000000000", 28068 => "0000000000000000", 28069 => "0000000000000000", 28070 => "0000000000000000", 28071 => "0000000000000000", 28072 => "0000000000000000", 28073 => "0000000000000000", 28074 => "0000000000000000", 28075 => "0000000000000000", 28076 => "0000000000000000", 28077 => "0000000000000000", 28078 => "0000000000000000", 28079 => "0000000000000000", 28080 => "0000000000000000", 28081 => "0000000000000000", 28082 => "0000000000000000", 28083 => "0000000000000000", 28084 => "0000000000000000", 28085 => "0000000000000000", 28086 => "0000000000000000", 28087 => "0000000000000000", 28088 => "0000000000000000", 28089 => "0000000000000000", 28090 => "0000000000000000", 28091 => "0000000000000000", 28092 => "0000000000000000", 28093 => "0000000000000000", 28094 => "0000000000000000", 28095 => "0000000000000000", 28096 => "0000000000000000", 28097 => "0000000000000000", 28098 => "0000000000000000", 28099 => "0000000000000000", 28100 => "0000000000000000", 28101 => "0000000000000000", 28102 => "0000000000000000", 28103 => "0000000000000000", 28104 => "0000000000000000", 28105 => "0000000000000000", 28106 => "0000000000000000", 28107 => "0000000000000000", 28108 => "0000000000000000", 28109 => "0000000000000000", 28110 => "0000000000000000", 28111 => "0000000000000000", 28112 => "0000000000000000", 28113 => "0000000000000000", 28114 => "0000000000000000", 28115 => "0000000000000000", 28116 => "0000000000000000", 28117 => "0000000000000000", 28118 => "0000000000000000", 28119 => "0000000000000000", 28120 => "0000000000000000", 28121 => "0000000000000000", 28122 => "0000000000000000", 28123 => "0000000000000000", 28124 => "0000000000000000", 28125 => "0000000000000000", 28126 => "0000000000000000", 28127 => "0000000000000000", 28128 => "0000000000000000", 28129 => "0000000000000000", 28130 => "0000000000000000", 28131 => "0000000000000000", 28132 => "0000000000000000", 28133 => "0000000000000000", 28134 => "0000000000000000", 28135 => "0000000000000000", 28136 => "0000000000000000", 28137 => "0000000000000000", 28138 => "0000000000000000", 28139 => "0000000000000000", 28140 => "0000000000000000", 28141 => "0000000000000000", 28142 => "0000000000000000", 28143 => "0000000000000000", 28144 => "0000000000000000", 28145 => "0000000000000000", 28146 => "0000000000000000", 28147 => "0000000000000000", 28148 => "0000000000000000", 28149 => "0000000000000000", 28150 => "0000000000000000", 28151 => "0000000000000000", 28152 => "0000000000000000", 28153 => "0000000000000000", 28154 => "0000000000000000", 28155 => "0000000000000000", 28156 => "0000000000000000", 28157 => "0000000000000000", 28158 => "0000000000000000", 28159 => "0000000000000000", 28160 => "0000000000000000", 28161 => "0000000000000000", 28162 => "0000000000000000", 28163 => "0000000000000000", 28164 => "0000000000000000", 28165 => "0000000000000000", 28166 => "0000000000000000", 28167 => "0000000000000000", 28168 => "0000000000000000", 28169 => "0000000000000000", 28170 => "0000000000000000", 28171 => "0000000000000000", 28172 => "0000000000000000", 28173 => "0000000000000000", 28174 => "0000000000000000", 28175 => "0000000000000000", 28176 => "0000000000000000", 28177 => "0000000000000000", 28178 => "0000000000000000", 28179 => "0000000000000000", 28180 => "0000000000000000", 28181 => "0000000000000000", 28182 => "0000000000000000", 28183 => "0000000000000000", 28184 => "0000000000000000", 28185 => "0000000000000000", 28186 => "0000000000000000", 28187 => "0000000000000000", 28188 => "0000000000000000", 28189 => "0000000000000000", 28190 => "0000000000000000", 28191 => "0000000000000000", 28192 => "0000000000000000", 28193 => "0000000000000000", 28194 => "0000000000000000", 28195 => "0000000000000000", 28196 => "0000000000000000", 28197 => "0000000000000000", 28198 => "0000000000000000", 28199 => "0000000000000000", 28200 => "0000000000000000", 28201 => "0000000000000000", 28202 => "0000000000000000", 28203 => "0000000000000000", 28204 => "0000000000000000", 28205 => "0000000000000000", 28206 => "0000000000000000", 28207 => "0000000000000000", 28208 => "0000000000000000", 28209 => "0000000000000000", 28210 => "0000000000000000", 28211 => "0000000000000000", 28212 => "0000000000000000", 28213 => "0000000000000000", 28214 => "0000000000000000", 28215 => "0000000000000000", 28216 => "0000000000000000", 28217 => "0000000000000000", 28218 => "0000000000000000", 28219 => "0000000000000000", 28220 => "0000000000000000", 28221 => "0000000000000000", 28222 => "0000000000000000", 28223 => "0000000000000000", 28224 => "0000000000000000", 28225 => "0000000000000000", 28226 => "0000000000000000", 28227 => "0000000000000000", 28228 => "0000000000000000", 28229 => "0000000000000000", 28230 => "0000000000000000", 28231 => "0000000000000000", 28232 => "0000000000000000", 28233 => "0000000000000000", 28234 => "0000000000000000", 28235 => "0000000000000000", 28236 => "0000000000000000", 28237 => "0000000000000000", 28238 => "0000000000000000", 28239 => "0000000000000000", 28240 => "0000000000000000", 28241 => "0000000000000000", 28242 => "0000000000000000", 28243 => "0000000000000000", 28244 => "0000000000000000", 28245 => "0000000000000000", 28246 => "0000000000000000", 28247 => "0000000000000000", 28248 => "0000000000000000", 28249 => "0000000000000000", 28250 => "0000000000000000", 28251 => "0000000000000000", 28252 => "0000000000000000", 28253 => "0000000000000000", 28254 => "0000000000000000", 28255 => "0000000000000000", 28256 => "0000000000000000", 28257 => "0000000000000000", 28258 => "0000000000000000", 28259 => "0000000000000000", 28260 => "0000000000000000", 28261 => "0000000000000000", 28262 => "0000000000000000", 28263 => "0000000000000000", 28264 => "0000000000000000", 28265 => "0000000000000000", 28266 => "0000000000000000", 28267 => "0000000000000000", 28268 => "0000000000000000", 28269 => "0000000000000000", 28270 => "0000000000000000", 28271 => "0000000000000000", 28272 => "0000000000000000", 28273 => "0000000000000000", 28274 => "0000000000000000", 28275 => "0000000000000000", 28276 => "0000000000000000", 28277 => "0000000000000000", 28278 => "0000000000000000", 28279 => "0000000000000000", 28280 => "0000000000000000", 28281 => "0000000000000000", 28282 => "0000000000000000", 28283 => "0000000000000000", 28284 => "0000000000000000", 28285 => "0000000000000000", 28286 => "0000000000000000", 28287 => "0000000000000000", 28288 => "0000000000000000", 28289 => "0000000000000000", 28290 => "0000000000000000", 28291 => "0000000000000000", 28292 => "0000000000000000", 28293 => "0000000000000000", 28294 => "0000000000000000", 28295 => "0000000000000000", 28296 => "0000000000000000", 28297 => "0000000000000000", 28298 => "0000000000000000", 28299 => "0000000000000000", 28300 => "0000000000000000", 28301 => "0000000000000000", 28302 => "0000000000000000", 28303 => "0000000000000000", 28304 => "0000000000000000", 28305 => "0000000000000000", 28306 => "0000000000000000", 28307 => "0000000000000000", 28308 => "0000000000000000", 28309 => "0000000000000000", 28310 => "0000000000000000", 28311 => "0000000000000000", 28312 => "0000000000000000", 28313 => "0000000000000000", 28314 => "0000000000000000", 28315 => "0000000000000000", 28316 => "0000000000000000", 28317 => "0000000000000000", 28318 => "0000000000000000", 28319 => "0000000000000000", 28320 => "0000000000000000", 28321 => "0000000000000000", 28322 => "0000000000000000", 28323 => "0000000000000000", 28324 => "0000000000000000", 28325 => "0000000000000000", 28326 => "0000000000000000", 28327 => "0000000000000000", 28328 => "0000000000000000", 28329 => "0000000000000000", 28330 => "0000000000000000", 28331 => "0000000000000000", 28332 => "0000000000000000", 28333 => "0000000000000000", 28334 => "0000000000000000", 28335 => "0000000000000000", 28336 => "0000000000000000", 28337 => "0000000000000000", 28338 => "0000000000000000", 28339 => "0000000000000000", 28340 => "0000000000000000", 28341 => "0000000000000000", 28342 => "0000000000000000", 28343 => "0000000000000000", 28344 => "0000000000000000", 28345 => "0000000000000000", 28346 => "0000000000000000", 28347 => "0000000000000000", 28348 => "0000000000000000", 28349 => "0000000000000000", 28350 => "0000000000000000", 28351 => "0000000000000000", 28352 => "0000000000000000", 28353 => "0000000000000000", 28354 => "0000000000000000", 28355 => "0000000000000000", 28356 => "0000000000000000", 28357 => "0000000000000000", 28358 => "0000000000000000", 28359 => "0000000000000000", 28360 => "0000000000000000", 28361 => "0000000000000000", 28362 => "0000000000000000", 28363 => "0000000000000000", 28364 => "0000000000000000", 28365 => "0000000000000000", 28366 => "0000000000000000", 28367 => "0000000000000000", 28368 => "0000000000000000", 28369 => "0000000000000000", 28370 => "0000000000000000", 28371 => "0000000000000000", 28372 => "0000000000000000", 28373 => "0000000000000000", 28374 => "0000000000000000", 28375 => "0000000000000000", 28376 => "0000000000000000", 28377 => "0000000000000000", 28378 => "0000000000000000", 28379 => "0000000000000000", 28380 => "0000000000000000", 28381 => "0000000000000000", 28382 => "0000000000000000", 28383 => "0000000000000000", 28384 => "0000000000000000", 28385 => "0000000000000000", 28386 => "0000000000000000", 28387 => "0000000000000000", 28388 => "0000000000000000", 28389 => "0000000000000000", 28390 => "0000000000000000", 28391 => "0000000000000000", 28392 => "0000000000000000", 28393 => "0000000000000000", 28394 => "0000000000000000", 28395 => "0000000000000000", 28396 => "0000000000000000", 28397 => "0000000000000000", 28398 => "0000000000000000", 28399 => "0000000000000000", 28400 => "0000000000000000", 28401 => "0000000000000000", 28402 => "0000000000000000", 28403 => "0000000000000000", 28404 => "0000000000000000", 28405 => "0000000000000000", 28406 => "0000000000000000", 28407 => "0000000000000000", 28408 => "0000000000000000", 28409 => "0000000000000000", 28410 => "0000000000000000", 28411 => "0000000000000000", 28412 => "0000000000000000", 28413 => "0000000000000000", 28414 => "0000000000000000", 28415 => "0000000000000000", 28416 => "0000000000000000", 28417 => "0000000000000000", 28418 => "0000000000000000", 28419 => "0000000000000000", 28420 => "0000000000000000", 28421 => "0000000000000000", 28422 => "0000000000000000", 28423 => "0000000000000000", 28424 => "0000000000000000", 28425 => "0000000000000000", 28426 => "0000000000000000", 28427 => "0000000000000000", 28428 => "0000000000000000", 28429 => "0000000000000000", 28430 => "0000000000000000", 28431 => "0000000000000000", 28432 => "0000000000000000", 28433 => "0000000000000000", 28434 => "0000000000000000", 28435 => "0000000000000000", 28436 => "0000000000000000", 28437 => "0000000000000000", 28438 => "0000000000000000", 28439 => "0000000000000000", 28440 => "0000000000000000", 28441 => "0000000000000000", 28442 => "0000000000000000", 28443 => "0000000000000000", 28444 => "0000000000000000", 28445 => "0000000000000000", 28446 => "0000000000000000", 28447 => "0000000000000000", 28448 => "0000000000000000", 28449 => "0000000000000000", 28450 => "0000000000000000", 28451 => "0000000000000000", 28452 => "0000000000000000", 28453 => "0000000000000000", 28454 => "0000000000000000", 28455 => "0000000000000000", 28456 => "0000000000000000", 28457 => "0000000000000000", 28458 => "0000000000000000", 28459 => "0000000000000000", 28460 => "0000000000000000", 28461 => "0000000000000000", 28462 => "0000000000000000", 28463 => "0000000000000000", 28464 => "0000000000000000", 28465 => "0000000000000000", 28466 => "0000000000000000", 28467 => "0000000000000000", 28468 => "0000000000000000", 28469 => "0000000000000000", 28470 => "0000000000000000", 28471 => "0000000000000000", 28472 => "0000000000000000", 28473 => "0000000000000000", 28474 => "0000000000000000", 28475 => "0000000000000000", 28476 => "0000000000000000", 28477 => "0000000000000000", 28478 => "0000000000000000", 28479 => "0000000000000000", 28480 => "0000000000000000", 28481 => "0000000000000000", 28482 => "0000000000000000", 28483 => "0000000000000000", 28484 => "0000000000000000", 28485 => "0000000000000000", 28486 => "0000000000000000", 28487 => "0000000000000000", 28488 => "0000000000000000", 28489 => "0000000000000000", 28490 => "0000000000000000", 28491 => "0000000000000000", 28492 => "0000000000000000", 28493 => "0000000000000000", 28494 => "0000000000000000", 28495 => "0000000000000000", 28496 => "0000000000000000", 28497 => "0000000000000000", 28498 => "0000000000000000", 28499 => "0000000000000000", 28500 => "0000000000000000", 28501 => "0000000000000000", 28502 => "0000000000000000", 28503 => "0000000000000000", 28504 => "0000000000000000", 28505 => "0000000000000000", 28506 => "0000000000000000", 28507 => "0000000000000000", 28508 => "0000000000000000", 28509 => "0000000000000000", 28510 => "0000000000000000", 28511 => "0000000000000000", 28512 => "0000000000000000", 28513 => "0000000000000000", 28514 => "0000000000000000", 28515 => "0000000000000000", 28516 => "0000000000000000", 28517 => "0000000000000000", 28518 => "0000000000000000", 28519 => "0000000000000000", 28520 => "0000000000000000", 28521 => "0000000000000000", 28522 => "0000000000000000", 28523 => "0000000000000000", 28524 => "0000000000000000", 28525 => "0000000000000000", 28526 => "0000000000000000", 28527 => "0000000000000000", 28528 => "0000000000000000", 28529 => "0000000000000000", 28530 => "0000000000000000", 28531 => "0000000000000000", 28532 => "0000000000000000", 28533 => "0000000000000000", 28534 => "0000000000000000", 28535 => "0000000000000000", 28536 => "0000000000000000", 28537 => "0000000000000000", 28538 => "0000000000000000", 28539 => "0000000000000000", 28540 => "0000000000000000", 28541 => "0000000000000000", 28542 => "0000000000000000", 28543 => "0000000000000000", 28544 => "0000000000000000", 28545 => "0000000000000000", 28546 => "0000000000000000", 28547 => "0000000000000000", 28548 => "0000000000000000", 28549 => "0000000000000000", 28550 => "0000000000000000", 28551 => "0000000000000000", 28552 => "0000000000000000", 28553 => "0000000000000000", 28554 => "0000000000000000", 28555 => "0000000000000000", 28556 => "0000000000000000", 28557 => "0000000000000000", 28558 => "0000000000000000", 28559 => "0000000000000000", 28560 => "0000000000000000", 28561 => "0000000000000000", 28562 => "0000000000000000", 28563 => "0000000000000000", 28564 => "0000000000000000", 28565 => "0000000000000000", 28566 => "0000000000000000", 28567 => "0000000000000000", 28568 => "0000000000000000", 28569 => "0000000000000000", 28570 => "0000000000000000", 28571 => "0000000000000000", 28572 => "0000000000000000", 28573 => "0000000000000000", 28574 => "0000000000000000", 28575 => "0000000000000000", 28576 => "0000000000000000", 28577 => "0000000000000000", 28578 => "0000000000000000", 28579 => "0000000000000000", 28580 => "0000000000000000", 28581 => "0000000000000000", 28582 => "0000000000000000", 28583 => "0000000000000000", 28584 => "0000000000000000", 28585 => "0000000000000000", 28586 => "0000000000000000", 28587 => "0000000000000000", 28588 => "0000000000000000", 28589 => "0000000000000000", 28590 => "0000000000000000", 28591 => "0000000000000000", 28592 => "0000000000000000", 28593 => "0000000000000000", 28594 => "0000000000000000", 28595 => "0000000000000000", 28596 => "0000000000000000", 28597 => "0000000000000000", 28598 => "0000000000000000", 28599 => "0000000000000000", 28600 => "0000000000000000", 28601 => "0000000000000000", 28602 => "0000000000000000", 28603 => "0000000000000000", 28604 => "0000000000000000", 28605 => "0000000000000000", 28606 => "0000000000000000", 28607 => "0000000000000000", 28608 => "0000000000000000", 28609 => "0000000000000000", 28610 => "0000000000000000", 28611 => "0000000000000000", 28612 => "0000000000000000", 28613 => "0000000000000000", 28614 => "0000000000000000", 28615 => "0000000000000000", 28616 => "0000000000000000", 28617 => "0000000000000000", 28618 => "0000000000000000", 28619 => "0000000000000000", 28620 => "0000000000000000", 28621 => "0000000000000000", 28622 => "0000000000000000", 28623 => "0000000000000000", 28624 => "0000000000000000", 28625 => "0000000000000000", 28626 => "0000000000000000", 28627 => "0000000000000000", 28628 => "0000000000000000", 28629 => "0000000000000000", 28630 => "0000000000000000", 28631 => "0000000000000000", 28632 => "0000000000000000", 28633 => "0000000000000000", 28634 => "0000000000000000", 28635 => "0000000000000000", 28636 => "0000000000000000", 28637 => "0000000000000000", 28638 => "0000000000000000", 28639 => "0000000000000000", 28640 => "0000000000000000", 28641 => "0000000000000000", 28642 => "0000000000000000", 28643 => "0000000000000000", 28644 => "0000000000000000", 28645 => "0000000000000000", 28646 => "0000000000000000", 28647 => "0000000000000000", 28648 => "0000000000000000", 28649 => "0000000000000000", 28650 => "0000000000000000", 28651 => "0000000000000000", 28652 => "0000000000000000", 28653 => "0000000000000000", 28654 => "0000000000000000", 28655 => "0000000000000000", 28656 => "0000000000000000", 28657 => "0000000000000000", 28658 => "0000000000000000", 28659 => "0000000000000000", 28660 => "0000000000000000", 28661 => "0000000000000000", 28662 => "0000000000000000", 28663 => "0000000000000000", 28664 => "0000000000000000", 28665 => "0000000000000000", 28666 => "0000000000000000", 28667 => "0000000000000000", 28668 => "0000000000000000", 28669 => "0000000000000000", 28670 => "0000000000000000", 28671 => "0000000000000000", 28672 => "0000000000000000", 28673 => "0000000000000000", 28674 => "0000000000000000", 28675 => "0000000000000000", 28676 => "0000000000000000", 28677 => "0000000000000000", 28678 => "0000000000000000", 28679 => "0000000000000000", 28680 => "0000000000000000", 28681 => "0000000000000000", 28682 => "0000000000000000", 28683 => "0000000000000000", 28684 => "0000000000000000", 28685 => "0000000000000000", 28686 => "0000000000000000", 28687 => "0000000000000000", 28688 => "0000000000000000", 28689 => "0000000000000000", 28690 => "0000000000000000", 28691 => "0000000000000000", 28692 => "0000000000000000", 28693 => "0000000000000000", 28694 => "0000000000000000", 28695 => "0000000000000000", 28696 => "0000000000000000", 28697 => "0000000000000000", 28698 => "0000000000000000", 28699 => "0000000000000000", 28700 => "0000000000000000", 28701 => "0000000000000000", 28702 => "0000000000000000", 28703 => "0000000000000000", 28704 => "0000000000000000", 28705 => "0000000000000000", 28706 => "0000000000000000", 28707 => "0000000000000000", 28708 => "0000000000000000", 28709 => "0000000000000000", 28710 => "0000000000000000", 28711 => "0000000000000000", 28712 => "0000000000000000", 28713 => "0000000000000000", 28714 => "0000000000000000", 28715 => "0000000000000000", 28716 => "0000000000000000", 28717 => "0000000000000000", 28718 => "0000000000000000", 28719 => "0000000000000000", 28720 => "0000000000000000", 28721 => "0000000000000000", 28722 => "0000000000000000", 28723 => "0000000000000000", 28724 => "0000000000000000", 28725 => "0000000000000000", 28726 => "0000000000000000", 28727 => "0000000000000000", 28728 => "0000000000000000", 28729 => "0000000000000000", 28730 => "0000000000000000", 28731 => "0000000000000000", 28732 => "0000000000000000", 28733 => "0000000000000000", 28734 => "0000000000000000", 28735 => "0000000000000000", 28736 => "0000000000000000", 28737 => "0000000000000000", 28738 => "0000000000000000", 28739 => "0000000000000000", 28740 => "0000000000000000", 28741 => "0000000000000000", 28742 => "0000000000000000", 28743 => "0000000000000000", 28744 => "0000000000000000", 28745 => "0000000000000000", 28746 => "0000000000000000", 28747 => "0000000000000000", 28748 => "0000000000000000", 28749 => "0000000000000000", 28750 => "0000000000000000", 28751 => "0000000000000000", 28752 => "0000000000000000", 28753 => "0000000000000000", 28754 => "0000000000000000", 28755 => "0000000000000000", 28756 => "0000000000000000", 28757 => "0000000000000000", 28758 => "0000000000000000", 28759 => "0000000000000000", 28760 => "0000000000000000", 28761 => "0000000000000000", 28762 => "0000000000000000", 28763 => "0000000000000000", 28764 => "0000000000000000", 28765 => "0000000000000000", 28766 => "0000000000000000", 28767 => "0000000000000000", 28768 => "0000000000000000", 28769 => "0000000000000000", 28770 => "0000000000000000", 28771 => "0000000000000000", 28772 => "0000000000000000", 28773 => "0000000000000000", 28774 => "0000000000000000", 28775 => "0000000000000000", 28776 => "0000000000000000", 28777 => "0000000000000000", 28778 => "0000000000000000", 28779 => "0000000000000000", 28780 => "0000000000000000", 28781 => "0000000000000000", 28782 => "0000000000000000", 28783 => "0000000000000000", 28784 => "0000000000000000", 28785 => "0000000000000000", 28786 => "0000000000000000", 28787 => "0000000000000000", 28788 => "0000000000000000", 28789 => "0000000000000000", 28790 => "0000000000000000", 28791 => "0000000000000000", 28792 => "0000000000000000", 28793 => "0000000000000000", 28794 => "0000000000000000", 28795 => "0000000000000000", 28796 => "0000000000000000", 28797 => "0000000000000000", 28798 => "0000000000000000", 28799 => "0000000000000000", 28800 => "0000000000000000", 28801 => "0000000000000000", 28802 => "0000000000000000", 28803 => "0000000000000000", 28804 => "0000000000000000", 28805 => "0000000000000000", 28806 => "0000000000000000", 28807 => "0000000000000000", 28808 => "0000000000000000", 28809 => "0000000000000000", 28810 => "0000000000000000", 28811 => "0000000000000000", 28812 => "0000000000000000", 28813 => "0000000000000000", 28814 => "0000000000000000", 28815 => "0000000000000000", 28816 => "0000000000000000", 28817 => "0000000000000000", 28818 => "0000000000000000", 28819 => "0000000000000000", 28820 => "0000000000000000", 28821 => "0000000000000000", 28822 => "0000000000000000", 28823 => "0000000000000000", 28824 => "0000000000000000", 28825 => "0000000000000000", 28826 => "0000000000000000", 28827 => "0000000000000000", 28828 => "0000000000000000", 28829 => "0000000000000000", 28830 => "0000000000000000", 28831 => "0000000000000000", 28832 => "0000000000000000", 28833 => "0000000000000000", 28834 => "0000000000000000", 28835 => "0000000000000000", 28836 => "0000000000000000", 28837 => "0000000000000000", 28838 => "0000000000000000", 28839 => "0000000000000000", 28840 => "0000000000000000", 28841 => "0000000000000000", 28842 => "0000000000000000", 28843 => "0000000000000000", 28844 => "0000000000000000", 28845 => "0000000000000000", 28846 => "0000000000000000", 28847 => "0000000000000000", 28848 => "0000000000000000", 28849 => "0000000000000000", 28850 => "0000000000000000", 28851 => "0000000000000000", 28852 => "0000000000000000", 28853 => "0000000000000000", 28854 => "0000000000000000", 28855 => "0000000000000000", 28856 => "0000000000000000", 28857 => "0000000000000000", 28858 => "0000000000000000", 28859 => "0000000000000000", 28860 => "0000000000000000", 28861 => "0000000000000000", 28862 => "0000000000000000", 28863 => "0000000000000000", 28864 => "0000000000000000", 28865 => "0000000000000000", 28866 => "0000000000000000", 28867 => "0000000000000000", 28868 => "0000000000000000", 28869 => "0000000000000000", 28870 => "0000000000000000", 28871 => "0000000000000000", 28872 => "0000000000000000", 28873 => "0000000000000000", 28874 => "0000000000000000", 28875 => "0000000000000000", 28876 => "0000000000000000", 28877 => "0000000000000000", 28878 => "0000000000000000", 28879 => "0000000000000000", 28880 => "0000000000000000", 28881 => "0000000000000000", 28882 => "0000000000000000", 28883 => "0000000000000000", 28884 => "0000000000000000", 28885 => "0000000000000000", 28886 => "0000000000000000", 28887 => "0000000000000000", 28888 => "0000000000000000", 28889 => "0000000000000000", 28890 => "0000000000000000", 28891 => "0000000000000000", 28892 => "0000000000000000", 28893 => "0000000000000000", 28894 => "0000000000000000", 28895 => "0000000000000000", 28896 => "0000000000000000", 28897 => "0000000000000000", 28898 => "0000000000000000", 28899 => "0000000000000000", 28900 => "0000000000000000", 28901 => "0000000000000000", 28902 => "0000000000000000", 28903 => "0000000000000000", 28904 => "0000000000000000", 28905 => "0000000000000000", 28906 => "0000000000000000", 28907 => "0000000000000000", 28908 => "0000000000000000", 28909 => "0000000000000000", 28910 => "0000000000000000", 28911 => "0000000000000000", 28912 => "0000000000000000", 28913 => "0000000000000000", 28914 => "0000000000000000", 28915 => "0000000000000000", 28916 => "0000000000000000", 28917 => "0000000000000000", 28918 => "0000000000000000", 28919 => "0000000000000000", 28920 => "0000000000000000", 28921 => "0000000000000000", 28922 => "0000000000000000", 28923 => "0000000000000000", 28924 => "0000000000000000", 28925 => "0000000000000000", 28926 => "0000000000000000", 28927 => "0000000000000000", 28928 => "0000000000000000", 28929 => "0000000000000000", 28930 => "0000000000000000", 28931 => "0000000000000000", 28932 => "0000000000000000", 28933 => "0000000000000000", 28934 => "0000000000000000", 28935 => "0000000000000000", 28936 => "0000000000000000", 28937 => "0000000000000000", 28938 => "0000000000000000", 28939 => "0000000000000000", 28940 => "0000000000000000", 28941 => "0000000000000000", 28942 => "0000000000000000", 28943 => "0000000000000000", 28944 => "0000000000000000", 28945 => "0000000000000000", 28946 => "0000000000000000", 28947 => "0000000000000000", 28948 => "0000000000000000", 28949 => "0000000000000000", 28950 => "0000000000000000", 28951 => "0000000000000000", 28952 => "0000000000000000", 28953 => "0000000000000000", 28954 => "0000000000000000", 28955 => "0000000000000000", 28956 => "0000000000000000", 28957 => "0000000000000000", 28958 => "0000000000000000", 28959 => "0000000000000000", 28960 => "0000000000000000", 28961 => "0000000000000000", 28962 => "0000000000000000", 28963 => "0000000000000000", 28964 => "0000000000000000", 28965 => "0000000000000000", 28966 => "0000000000000000", 28967 => "0000000000000000", 28968 => "0000000000000000", 28969 => "0000000000000000", 28970 => "0000000000000000", 28971 => "0000000000000000", 28972 => "0000000000000000", 28973 => "0000000000000000", 28974 => "0000000000000000", 28975 => "0000000000000000", 28976 => "0000000000000000", 28977 => "0000000000000000", 28978 => "0000000000000000", 28979 => "0000000000000000", 28980 => "0000000000000000", 28981 => "0000000000000000", 28982 => "0000000000000000", 28983 => "0000000000000000", 28984 => "0000000000000000", 28985 => "0000000000000000", 28986 => "0000000000000000", 28987 => "0000000000000000", 28988 => "0000000000000000", 28989 => "0000000000000000", 28990 => "0000000000000000", 28991 => "0000000000000000", 28992 => "0000000000000000", 28993 => "0000000000000000", 28994 => "0000000000000000", 28995 => "0000000000000000", 28996 => "0000000000000000", 28997 => "0000000000000000", 28998 => "0000000000000000", 28999 => "0000000000000000", 29000 => "0000000000000000", 29001 => "0000000000000000", 29002 => "0000000000000000", 29003 => "0000000000000000", 29004 => "0000000000000000", 29005 => "0000000000000000", 29006 => "0000000000000000", 29007 => "0000000000000000", 29008 => "0000000000000000", 29009 => "0000000000000000", 29010 => "0000000000000000", 29011 => "0000000000000000", 29012 => "0000000000000000", 29013 => "0000000000000000", 29014 => "0000000000000000", 29015 => "0000000000000000", 29016 => "0000000000000000", 29017 => "0000000000000000", 29018 => "0000000000000000", 29019 => "0000000000000000", 29020 => "0000000000000000", 29021 => "0000000000000000", 29022 => "0000000000000000", 29023 => "0000000000000000", 29024 => "0000000000000000", 29025 => "0000000000000000", 29026 => "0000000000000000", 29027 => "0000000000000000", 29028 => "0000000000000000", 29029 => "0000000000000000", 29030 => "0000000000000000", 29031 => "0000000000000000", 29032 => "0000000000000000", 29033 => "0000000000000000", 29034 => "0000000000000000", 29035 => "0000000000000000", 29036 => "0000000000000000", 29037 => "0000000000000000", 29038 => "0000000000000000", 29039 => "0000000000000000", 29040 => "0000000000000000", 29041 => "0000000000000000", 29042 => "0000000000000000", 29043 => "0000000000000000", 29044 => "0000000000000000", 29045 => "0000000000000000", 29046 => "0000000000000000", 29047 => "0000000000000000", 29048 => "0000000000000000", 29049 => "0000000000000000", 29050 => "0000000000000000", 29051 => "0000000000000000", 29052 => "0000000000000000", 29053 => "0000000000000000", 29054 => "0000000000000000", 29055 => "0000000000000000", 29056 => "0000000000000000", 29057 => "0000000000000000", 29058 => "0000000000000000", 29059 => "0000000000000000", 29060 => "0000000000000000", 29061 => "0000000000000000", 29062 => "0000000000000000", 29063 => "0000000000000000", 29064 => "0000000000000000", 29065 => "0000000000000000", 29066 => "0000000000000000", 29067 => "0000000000000000", 29068 => "0000000000000000", 29069 => "0000000000000000", 29070 => "0000000000000000", 29071 => "0000000000000000", 29072 => "0000000000000000", 29073 => "0000000000000000", 29074 => "0000000000000000", 29075 => "0000000000000000", 29076 => "0000000000000000", 29077 => "0000000000000000", 29078 => "0000000000000000", 29079 => "0000000000000000", 29080 => "0000000000000000", 29081 => "0000000000000000", 29082 => "0000000000000000", 29083 => "0000000000000000", 29084 => "0000000000000000", 29085 => "0000000000000000", 29086 => "0000000000000000", 29087 => "0000000000000000", 29088 => "0000000000000000", 29089 => "0000000000000000", 29090 => "0000000000000000", 29091 => "0000000000000000", 29092 => "0000000000000000", 29093 => "0000000000000000", 29094 => "0000000000000000", 29095 => "0000000000000000", 29096 => "0000000000000000", 29097 => "0000000000000000", 29098 => "0000000000000000", 29099 => "0000000000000000", 29100 => "0000000000000000", 29101 => "0000000000000000", 29102 => "0000000000000000", 29103 => "0000000000000000", 29104 => "0000000000000000", 29105 => "0000000000000000", 29106 => "0000000000000000", 29107 => "0000000000000000", 29108 => "0000000000000000", 29109 => "0000000000000000", 29110 => "0000000000000000", 29111 => "0000000000000000", 29112 => "0000000000000000", 29113 => "0000000000000000", 29114 => "0000000000000000", 29115 => "0000000000000000", 29116 => "0000000000000000", 29117 => "0000000000000000", 29118 => "0000000000000000", 29119 => "0000000000000000", 29120 => "0000000000000000", 29121 => "0000000000000000", 29122 => "0000000000000000", 29123 => "0000000000000000", 29124 => "0000000000000000", 29125 => "0000000000000000", 29126 => "0000000000000000", 29127 => "0000000000000000", 29128 => "0000000000000000", 29129 => "0000000000000000", 29130 => "0000000000000000", 29131 => "0000000000000000", 29132 => "0000000000000000", 29133 => "0000000000000000", 29134 => "0000000000000000", 29135 => "0000000000000000", 29136 => "0000000000000000", 29137 => "0000000000000000", 29138 => "0000000000000000", 29139 => "0000000000000000", 29140 => "0000000000000000", 29141 => "0000000000000000", 29142 => "0000000000000000", 29143 => "0000000000000000", 29144 => "0000000000000000", 29145 => "0000000000000000", 29146 => "0000000000000000", 29147 => "0000000000000000", 29148 => "0000000000000000", 29149 => "0000000000000000", 29150 => "0000000000000000", 29151 => "0000000000000000", 29152 => "0000000000000000", 29153 => "0000000000000000", 29154 => "0000000000000000", 29155 => "0000000000000000", 29156 => "0000000000000000", 29157 => "0000000000000000", 29158 => "0000000000000000", 29159 => "0000000000000000", 29160 => "0000000000000000", 29161 => "0000000000000000", 29162 => "0000000000000000", 29163 => "0000000000000000", 29164 => "0000000000000000", 29165 => "0000000000000000", 29166 => "0000000000000000", 29167 => "0000000000000000", 29168 => "0000000000000000", 29169 => "0000000000000000", 29170 => "0000000000000000", 29171 => "0000000000000000", 29172 => "0000000000000000", 29173 => "0000000000000000", 29174 => "0000000000000000", 29175 => "0000000000000000", 29176 => "0000000000000000", 29177 => "0000000000000000", 29178 => "0000000000000000", 29179 => "0000000000000000", 29180 => "0000000000000000", 29181 => "0000000000000000", 29182 => "0000000000000000", 29183 => "0000000000000000", 29184 => "0000000000000000", 29185 => "0000000000000000", 29186 => "0000000000000000", 29187 => "0000000000000000", 29188 => "0000000000000000", 29189 => "0000000000000000", 29190 => "0000000000000000", 29191 => "0000000000000000", 29192 => "0000000000000000", 29193 => "0000000000000000", 29194 => "0000000000000000", 29195 => "0000000000000000", 29196 => "0000000000000000", 29197 => "0000000000000000", 29198 => "0000000000000000", 29199 => "0000000000000000", 29200 => "0000000000000000", 29201 => "0000000000000000", 29202 => "0000000000000000", 29203 => "0000000000000000", 29204 => "0000000000000000", 29205 => "0000000000000000", 29206 => "0000000000000000", 29207 => "0000000000000000", 29208 => "0000000000000000", 29209 => "0000000000000000", 29210 => "0000000000000000", 29211 => "0000000000000000", 29212 => "0000000000000000", 29213 => "0000000000000000", 29214 => "0000000000000000", 29215 => "0000000000000000", 29216 => "0000000000000000", 29217 => "0000000000000000", 29218 => "0000000000000000", 29219 => "0000000000000000", 29220 => "0000000000000000", 29221 => "0000000000000000", 29222 => "0000000000000000", 29223 => "0000000000000000", 29224 => "0000000000000000", 29225 => "0000000000000000", 29226 => "0000000000000000", 29227 => "0000000000000000", 29228 => "0000000000000000", 29229 => "0000000000000000", 29230 => "0000000000000000", 29231 => "0000000000000000", 29232 => "0000000000000000", 29233 => "0000000000000000", 29234 => "0000000000000000", 29235 => "0000000000000000", 29236 => "0000000000000000", 29237 => "0000000000000000", 29238 => "0000000000000000", 29239 => "0000000000000000", 29240 => "0000000000000000", 29241 => "0000000000000000", 29242 => "0000000000000000", 29243 => "0000000000000000", 29244 => "0000000000000000", 29245 => "0000000000000000", 29246 => "0000000000000000", 29247 => "0000000000000000", 29248 => "0000000000000000", 29249 => "0000000000000000", 29250 => "0000000000000000", 29251 => "0000000000000000", 29252 => "0000000000000000", 29253 => "0000000000000000", 29254 => "0000000000000000", 29255 => "0000000000000000", 29256 => "0000000000000000", 29257 => "0000000000000000", 29258 => "0000000000000000", 29259 => "0000000000000000", 29260 => "0000000000000000", 29261 => "0000000000000000", 29262 => "0000000000000000", 29263 => "0000000000000000", 29264 => "0000000000000000", 29265 => "0000000000000000", 29266 => "0000000000000000", 29267 => "0000000000000000", 29268 => "0000000000000000", 29269 => "0000000000000000", 29270 => "0000000000000000", 29271 => "0000000000000000", 29272 => "0000000000000000", 29273 => "0000000000000000", 29274 => "0000000000000000", 29275 => "0000000000000000", 29276 => "0000000000000000", 29277 => "0000000000000000", 29278 => "0000000000000000", 29279 => "0000000000000000", 29280 => "0000000000000000", 29281 => "0000000000000000", 29282 => "0000000000000000", 29283 => "0000000000000000", 29284 => "0000000000000000", 29285 => "0000000000000000", 29286 => "0000000000000000", 29287 => "0000000000000000", 29288 => "0000000000000000", 29289 => "0000000000000000", 29290 => "0000000000000000", 29291 => "0000000000000000", 29292 => "0000000000000000", 29293 => "0000000000000000", 29294 => "0000000000000000", 29295 => "0000000000000000", 29296 => "0000000000000000", 29297 => "0000000000000000", 29298 => "0000000000000000", 29299 => "0000000000000000", 29300 => "0000000000000000", 29301 => "0000000000000000", 29302 => "0000000000000000", 29303 => "0000000000000000", 29304 => "0000000000000000", 29305 => "0000000000000000", 29306 => "0000000000000000", 29307 => "0000000000000000", 29308 => "0000000000000000", 29309 => "0000000000000000", 29310 => "0000000000000000", 29311 => "0000000000000000", 29312 => "0000000000000000", 29313 => "0000000000000000", 29314 => "0000000000000000", 29315 => "0000000000000000", 29316 => "0000000000000000", 29317 => "0000000000000000", 29318 => "0000000000000000", 29319 => "0000000000000000", 29320 => "0000000000000000", 29321 => "0000000000000000", 29322 => "0000000000000000", 29323 => "0000000000000000", 29324 => "0000000000000000", 29325 => "0000000000000000", 29326 => "0000000000000000", 29327 => "0000000000000000", 29328 => "0000000000000000", 29329 => "0000000000000000", 29330 => "0000000000000000", 29331 => "0000000000000000", 29332 => "0000000000000000", 29333 => "0000000000000000", 29334 => "0000000000000000", 29335 => "0000000000000000", 29336 => "0000000000000000", 29337 => "0000000000000000", 29338 => "0000000000000000", 29339 => "0000000000000000", 29340 => "0000000000000000", 29341 => "0000000000000000", 29342 => "0000000000000000", 29343 => "0000000000000000", 29344 => "0000000000000000", 29345 => "0000000000000000", 29346 => "0000000000000000", 29347 => "0000000000000000", 29348 => "0000000000000000", 29349 => "0000000000000000", 29350 => "0000000000000000", 29351 => "0000000000000000", 29352 => "0000000000000000", 29353 => "0000000000000000", 29354 => "0000000000000000", 29355 => "0000000000000000", 29356 => "0000000000000000", 29357 => "0000000000000000", 29358 => "0000000000000000", 29359 => "0000000000000000", 29360 => "0000000000000000", 29361 => "0000000000000000", 29362 => "0000000000000000", 29363 => "0000000000000000", 29364 => "0000000000000000", 29365 => "0000000000000000", 29366 => "0000000000000000", 29367 => "0000000000000000", 29368 => "0000000000000000", 29369 => "0000000000000000", 29370 => "0000000000000000", 29371 => "0000000000000000", 29372 => "0000000000000000", 29373 => "0000000000000000", 29374 => "0000000000000000", 29375 => "0000000000000000", 29376 => "0000000000000000", 29377 => "0000000000000000", 29378 => "0000000000000000", 29379 => "0000000000000000", 29380 => "0000000000000000", 29381 => "0000000000000000", 29382 => "0000000000000000", 29383 => "0000000000000000", 29384 => "0000000000000000", 29385 => "0000000000000000", 29386 => "0000000000000000", 29387 => "0000000000000000", 29388 => "0000000000000000", 29389 => "0000000000000000", 29390 => "0000000000000000", 29391 => "0000000000000000", 29392 => "0000000000000000", 29393 => "0000000000000000", 29394 => "0000000000000000", 29395 => "0000000000000000", 29396 => "0000000000000000", 29397 => "0000000000000000", 29398 => "0000000000000000", 29399 => "0000000000000000", 29400 => "0000000000000000", 29401 => "0000000000000000", 29402 => "0000000000000000", 29403 => "0000000000000000", 29404 => "0000000000000000", 29405 => "0000000000000000", 29406 => "0000000000000000", 29407 => "0000000000000000", 29408 => "0000000000000000", 29409 => "0000000000000000", 29410 => "0000000000000000", 29411 => "0000000000000000", 29412 => "0000000000000000", 29413 => "0000000000000000", 29414 => "0000000000000000", 29415 => "0000000000000000", 29416 => "0000000000000000", 29417 => "0000000000000000", 29418 => "0000000000000000", 29419 => "0000000000000000", 29420 => "0000000000000000", 29421 => "0000000000000000", 29422 => "0000000000000000", 29423 => "0000000000000000", 29424 => "0000000000000000", 29425 => "0000000000000000", 29426 => "0000000000000000", 29427 => "0000000000000000", 29428 => "0000000000000000", 29429 => "0000000000000000", 29430 => "0000000000000000", 29431 => "0000000000000000", 29432 => "0000000000000000", 29433 => "0000000000000000", 29434 => "0000000000000000", 29435 => "0000000000000000", 29436 => "0000000000000000", 29437 => "0000000000000000", 29438 => "0000000000000000", 29439 => "0000000000000000", 29440 => "0000000000000000", 29441 => "0000000000000000", 29442 => "0000000000000000", 29443 => "0000000000000000", 29444 => "0000000000000000", 29445 => "0000000000000000", 29446 => "0000000000000000", 29447 => "0000000000000000", 29448 => "0000000000000000", 29449 => "0000000000000000", 29450 => "0000000000000000", 29451 => "0000000000000000", 29452 => "0000000000000000", 29453 => "0000000000000000", 29454 => "0000000000000000", 29455 => "0000000000000000", 29456 => "0000000000000000", 29457 => "0000000000000000", 29458 => "0000000000000000", 29459 => "0000000000000000", 29460 => "0000000000000000", 29461 => "0000000000000000", 29462 => "0000000000000000", 29463 => "0000000000000000", 29464 => "0000000000000000", 29465 => "0000000000000000", 29466 => "0000000000000000", 29467 => "0000000000000000", 29468 => "0000000000000000", 29469 => "0000000000000000", 29470 => "0000000000000000", 29471 => "0000000000000000", 29472 => "0000000000000000", 29473 => "0000000000000000", 29474 => "0000000000000000", 29475 => "0000000000000000", 29476 => "0000000000000000", 29477 => "0000000000000000", 29478 => "0000000000000000", 29479 => "0000000000000000", 29480 => "0000000000000000", 29481 => "0000000000000000", 29482 => "0000000000000000", 29483 => "0000000000000000", 29484 => "0000000000000000", 29485 => "0000000000000000", 29486 => "0000000000000000", 29487 => "0000000000000000", 29488 => "0000000000000000", 29489 => "0000000000000000", 29490 => "0000000000000000", 29491 => "0000000000000000", 29492 => "0000000000000000", 29493 => "0000000000000000", 29494 => "0000000000000000", 29495 => "0000000000000000", 29496 => "0000000000000000", 29497 => "0000000000000000", 29498 => "0000000000000000", 29499 => "0000000000000000", 29500 => "0000000000000000", 29501 => "0000000000000000", 29502 => "0000000000000000", 29503 => "0000000000000000", 29504 => "0000000000000000", 29505 => "0000000000000000", 29506 => "0000000000000000", 29507 => "0000000000000000", 29508 => "0000000000000000", 29509 => "0000000000000000", 29510 => "0000000000000000", 29511 => "0000000000000000", 29512 => "0000000000000000", 29513 => "0000000000000000", 29514 => "0000000000000000", 29515 => "0000000000000000", 29516 => "0000000000000000", 29517 => "0000000000000000", 29518 => "0000000000000000", 29519 => "0000000000000000", 29520 => "0000000000000000", 29521 => "0000000000000000", 29522 => "0000000000000000", 29523 => "0000000000000000", 29524 => "0000000000000000", 29525 => "0000000000000000", 29526 => "0000000000000000", 29527 => "0000000000000000", 29528 => "0000000000000000", 29529 => "0000000000000000", 29530 => "0000000000000000", 29531 => "0000000000000000", 29532 => "0000000000000000", 29533 => "0000000000000000", 29534 => "0000000000000000", 29535 => "0000000000000000", 29536 => "0000000000000000", 29537 => "0000000000000000", 29538 => "0000000000000000", 29539 => "0000000000000000", 29540 => "0000000000000000", 29541 => "0000000000000000", 29542 => "0000000000000000", 29543 => "0000000000000000", 29544 => "0000000000000000", 29545 => "0000000000000000", 29546 => "0000000000000000", 29547 => "0000000000000000", 29548 => "0000000000000000", 29549 => "0000000000000000", 29550 => "0000000000000000", 29551 => "0000000000000000", 29552 => "0000000000000000", 29553 => "0000000000000000", 29554 => "0000000000000000", 29555 => "0000000000000000", 29556 => "0000000000000000", 29557 => "0000000000000000", 29558 => "0000000000000000", 29559 => "0000000000000000", 29560 => "0000000000000000", 29561 => "0000000000000000", 29562 => "0000000000000000", 29563 => "0000000000000000", 29564 => "0000000000000000", 29565 => "0000000000000000", 29566 => "0000000000000000", 29567 => "0000000000000000", 29568 => "0000000000000000", 29569 => "0000000000000000", 29570 => "0000000000000000", 29571 => "0000000000000000", 29572 => "0000000000000000", 29573 => "0000000000000000", 29574 => "0000000000000000", 29575 => "0000000000000000", 29576 => "0000000000000000", 29577 => "0000000000000000", 29578 => "0000000000000000", 29579 => "0000000000000000", 29580 => "0000000000000000", 29581 => "0000000000000000", 29582 => "0000000000000000", 29583 => "0000000000000000", 29584 => "0000000000000000", 29585 => "0000000000000000", 29586 => "0000000000000000", 29587 => "0000000000000000", 29588 => "0000000000000000", 29589 => "0000000000000000", 29590 => "0000000000000000", 29591 => "0000000000000000", 29592 => "0000000000000000", 29593 => "0000000000000000", 29594 => "0000000000000000", 29595 => "0000000000000000", 29596 => "0000000000000000", 29597 => "0000000000000000", 29598 => "0000000000000000", 29599 => "0000000000000000", 29600 => "0000000000000000", 29601 => "0000000000000000", 29602 => "0000000000000000", 29603 => "0000000000000000", 29604 => "0000000000000000", 29605 => "0000000000000000", 29606 => "0000000000000000", 29607 => "0000000000000000", 29608 => "0000000000000000", 29609 => "0000000000000000", 29610 => "0000000000000000", 29611 => "0000000000000000", 29612 => "0000000000000000", 29613 => "0000000000000000", 29614 => "0000000000000000", 29615 => "0000000000000000", 29616 => "0000000000000000", 29617 => "0000000000000000", 29618 => "0000000000000000", 29619 => "0000000000000000", 29620 => "0000000000000000", 29621 => "0000000000000000", 29622 => "0000000000000000", 29623 => "0000000000000000", 29624 => "0000000000000000", 29625 => "0000000000000000", 29626 => "0000000000000000", 29627 => "0000000000000000", 29628 => "0000000000000000", 29629 => "0000000000000000", 29630 => "0000000000000000", 29631 => "0000000000000000", 29632 => "0000000000000000", 29633 => "0000000000000000", 29634 => "0000000000000000", 29635 => "0000000000000000", 29636 => "0000000000000000", 29637 => "0000000000000000", 29638 => "0000000000000000", 29639 => "0000000000000000", 29640 => "0000000000000000", 29641 => "0000000000000000", 29642 => "0000000000000000", 29643 => "0000000000000000", 29644 => "0000000000000000", 29645 => "0000000000000000", 29646 => "0000000000000000", 29647 => "0000000000000000", 29648 => "0000000000000000", 29649 => "0000000000000000", 29650 => "0000000000000000", 29651 => "0000000000000000", 29652 => "0000000000000000", 29653 => "0000000000000000", 29654 => "0000000000000000", 29655 => "0000000000000000", 29656 => "0000000000000000", 29657 => "0000000000000000", 29658 => "0000000000000000", 29659 => "0000000000000000", 29660 => "0000000000000000", 29661 => "0000000000000000", 29662 => "0000000000000000", 29663 => "0000000000000000", 29664 => "0000000000000000", 29665 => "0000000000000000", 29666 => "0000000000000000", 29667 => "0000000000000000", 29668 => "0000000000000000", 29669 => "0000000000000000", 29670 => "0000000000000000", 29671 => "0000000000000000", 29672 => "0000000000000000", 29673 => "0000000000000000", 29674 => "0000000000000000", 29675 => "0000000000000000", 29676 => "0000000000000000", 29677 => "0000000000000000", 29678 => "0000000000000000", 29679 => "0000000000000000", 29680 => "0000000000000000", 29681 => "0000000000000000", 29682 => "0000000000000000", 29683 => "0000000000000000", 29684 => "0000000000000000", 29685 => "0000000000000000", 29686 => "0000000000000000", 29687 => "0000000000000000", 29688 => "0000000000000000", 29689 => "0000000000000000", 29690 => "0000000000000000", 29691 => "0000000000000000", 29692 => "0000000000000000", 29693 => "0000000000000000", 29694 => "0000000000000000", 29695 => "0000000000000000", 29696 => "0000000000000000", 29697 => "0000000000000000", 29698 => "0000000000000000", 29699 => "0000000000000000", 29700 => "0000000000000000", 29701 => "0000000000000000", 29702 => "0000000000000000", 29703 => "0000000000000000", 29704 => "0000000000000000", 29705 => "0000000000000000", 29706 => "0000000000000000", 29707 => "0000000000000000", 29708 => "0000000000000000", 29709 => "0000000000000000", 29710 => "0000000000000000", 29711 => "0000000000000000", 29712 => "0000000000000000", 29713 => "0000000000000000", 29714 => "0000000000000000", 29715 => "0000000000000000", 29716 => "0000000000000000", 29717 => "0000000000000000", 29718 => "0000000000000000", 29719 => "0000000000000000", 29720 => "0000000000000000", 29721 => "0000000000000000", 29722 => "0000000000000000", 29723 => "0000000000000000", 29724 => "0000000000000000", 29725 => "0000000000000000", 29726 => "0000000000000000", 29727 => "0000000000000000", 29728 => "0000000000000000", 29729 => "0000000000000000", 29730 => "0000000000000000", 29731 => "0000000000000000", 29732 => "0000000000000000", 29733 => "0000000000000000", 29734 => "0000000000000000", 29735 => "0000000000000000", 29736 => "0000000000000000", 29737 => "0000000000000000", 29738 => "0000000000000000", 29739 => "0000000000000000", 29740 => "0000000000000000", 29741 => "0000000000000000", 29742 => "0000000000000000", 29743 => "0000000000000000", 29744 => "0000000000000000", 29745 => "0000000000000000", 29746 => "0000000000000000", 29747 => "0000000000000000", 29748 => "0000000000000000", 29749 => "0000000000000000", 29750 => "0000000000000000", 29751 => "0000000000000000", 29752 => "0000000000000000", 29753 => "0000000000000000", 29754 => "0000000000000000", 29755 => "0000000000000000", 29756 => "0000000000000000", 29757 => "0000000000000000", 29758 => "0000000000000000", 29759 => "0000000000000000", 29760 => "0000000000000000", 29761 => "0000000000000000", 29762 => "0000000000000000", 29763 => "0000000000000000", 29764 => "0000000000000000", 29765 => "0000000000000000", 29766 => "0000000000000000", 29767 => "0000000000000000", 29768 => "0000000000000000", 29769 => "0000000000000000", 29770 => "0000000000000000", 29771 => "0000000000000000", 29772 => "0000000000000000", 29773 => "0000000000000000", 29774 => "0000000000000000", 29775 => "0000000000000000", 29776 => "0000000000000000", 29777 => "0000000000000000", 29778 => "0000000000000000", 29779 => "0000000000000000", 29780 => "0000000000000000", 29781 => "0000000000000000", 29782 => "0000000000000000", 29783 => "0000000000000000", 29784 => "0000000000000000", 29785 => "0000000000000000", 29786 => "0000000000000000", 29787 => "0000000000000000", 29788 => "0000000000000000", 29789 => "0000000000000000", 29790 => "0000000000000000", 29791 => "0000000000000000", 29792 => "0000000000000000", 29793 => "0000000000000000", 29794 => "0000000000000000", 29795 => "0000000000000000", 29796 => "0000000000000000", 29797 => "0000000000000000", 29798 => "0000000000000000", 29799 => "0000000000000000", 29800 => "0000000000000000", 29801 => "0000000000000000", 29802 => "0000000000000000", 29803 => "0000000000000000", 29804 => "0000000000000000", 29805 => "0000000000000000", 29806 => "0000000000000000", 29807 => "0000000000000000", 29808 => "0000000000000000", 29809 => "0000000000000000", 29810 => "0000000000000000", 29811 => "0000000000000000", 29812 => "0000000000000000", 29813 => "0000000000000000", 29814 => "0000000000000000", 29815 => "0000000000000000", 29816 => "0000000000000000", 29817 => "0000000000000000", 29818 => "0000000000000000", 29819 => "0000000000000000", 29820 => "0000000000000000", 29821 => "0000000000000000", 29822 => "0000000000000000", 29823 => "0000000000000000", 29824 => "0000000000000000", 29825 => "0000000000000000", 29826 => "0000000000000000", 29827 => "0000000000000000", 29828 => "0000000000000000", 29829 => "0000000000000000", 29830 => "0000000000000000", 29831 => "0000000000000000", 29832 => "0000000000000000", 29833 => "0000000000000000", 29834 => "0000000000000000", 29835 => "0000000000000000", 29836 => "0000000000000000", 29837 => "0000000000000000", 29838 => "0000000000000000", 29839 => "0000000000000000", 29840 => "0000000000000000", 29841 => "0000000000000000", 29842 => "0000000000000000", 29843 => "0000000000000000", 29844 => "0000000000000000", 29845 => "0000000000000000", 29846 => "0000000000000000", 29847 => "0000000000000000", 29848 => "0000000000000000", 29849 => "0000000000000000", 29850 => "0000000000000000", 29851 => "0000000000000000", 29852 => "0000000000000000", 29853 => "0000000000000000", 29854 => "0000000000000000", 29855 => "0000000000000000", 29856 => "0000000000000000", 29857 => "0000000000000000", 29858 => "0000000000000000", 29859 => "0000000000000000", 29860 => "0000000000000000", 29861 => "0000000000000000", 29862 => "0000000000000000", 29863 => "0000000000000000", 29864 => "0000000000000000", 29865 => "0000000000000000", 29866 => "0000000000000000", 29867 => "0000000000000000", 29868 => "0000000000000000", 29869 => "0000000000000000", 29870 => "0000000000000000", 29871 => "0000000000000000", 29872 => "0000000000000000", 29873 => "0000000000000000", 29874 => "0000000000000000", 29875 => "0000000000000000", 29876 => "0000000000000000", 29877 => "0000000000000000", 29878 => "0000000000000000", 29879 => "0000000000000000", 29880 => "0000000000000000", 29881 => "0000000000000000", 29882 => "0000000000000000", 29883 => "0000000000000000", 29884 => "0000000000000000", 29885 => "0000000000000000", 29886 => "0000000000000000", 29887 => "0000000000000000", 29888 => "0000000000000000", 29889 => "0000000000000000", 29890 => "0000000000000000", 29891 => "0000000000000000", 29892 => "0000000000000000", 29893 => "0000000000000000", 29894 => "0000000000000000", 29895 => "0000000000000000", 29896 => "0000000000000000", 29897 => "0000000000000000", 29898 => "0000000000000000", 29899 => "0000000000000000", 29900 => "0000000000000000", 29901 => "0000000000000000", 29902 => "0000000000000000", 29903 => "0000000000000000", 29904 => "0000000000000000", 29905 => "0000000000000000", 29906 => "0000000000000000", 29907 => "0000000000000000", 29908 => "0000000000000000", 29909 => "0000000000000000", 29910 => "0000000000000000", 29911 => "0000000000000000", 29912 => "0000000000000000", 29913 => "0000000000000000", 29914 => "0000000000000000", 29915 => "0000000000000000", 29916 => "0000000000000000", 29917 => "0000000000000000", 29918 => "0000000000000000", 29919 => "0000000000000000", 29920 => "0000000000000000", 29921 => "0000000000000000", 29922 => "0000000000000000", 29923 => "0000000000000000", 29924 => "0000000000000000", 29925 => "0000000000000000", 29926 => "0000000000000000", 29927 => "0000000000000000", 29928 => "0000000000000000", 29929 => "0000000000000000", 29930 => "0000000000000000", 29931 => "0000000000000000", 29932 => "0000000000000000", 29933 => "0000000000000000", 29934 => "0000000000000000", 29935 => "0000000000000000", 29936 => "0000000000000000", 29937 => "0000000000000000", 29938 => "0000000000000000", 29939 => "0000000000000000", 29940 => "0000000000000000", 29941 => "0000000000000000", 29942 => "0000000000000000", 29943 => "0000000000000000", 29944 => "0000000000000000", 29945 => "0000000000000000", 29946 => "0000000000000000", 29947 => "0000000000000000", 29948 => "0000000000000000", 29949 => "0000000000000000", 29950 => "0000000000000000", 29951 => "0000000000000000", 29952 => "0000000000000000", 29953 => "0000000000000000", 29954 => "0000000000000000", 29955 => "0000000000000000", 29956 => "0000000000000000", 29957 => "0000000000000000", 29958 => "0000000000000000", 29959 => "0000000000000000", 29960 => "0000000000000000", 29961 => "0000000000000000", 29962 => "0000000000000000", 29963 => "0000000000000000", 29964 => "0000000000000000", 29965 => "0000000000000000", 29966 => "0000000000000000", 29967 => "0000000000000000", 29968 => "0000000000000000", 29969 => "0000000000000000", 29970 => "0000000000000000", 29971 => "0000000000000000", 29972 => "0000000000000000", 29973 => "0000000000000000", 29974 => "0000000000000000", 29975 => "0000000000000000", 29976 => "0000000000000000", 29977 => "0000000000000000", 29978 => "0000000000000000", 29979 => "0000000000000000", 29980 => "0000000000000000", 29981 => "0000000000000000", 29982 => "0000000000000000", 29983 => "0000000000000000", 29984 => "0000000000000000", 29985 => "0000000000000000", 29986 => "0000000000000000", 29987 => "0000000000000000", 29988 => "0000000000000000", 29989 => "0000000000000000", 29990 => "0000000000000000", 29991 => "0000000000000000", 29992 => "0000000000000000", 29993 => "0000000000000000", 29994 => "0000000000000000", 29995 => "0000000000000000", 29996 => "0000000000000000", 29997 => "0000000000000000", 29998 => "0000000000000000", 29999 => "0000000000000000", 30000 => "0000000000000000", 30001 => "0000000000000000", 30002 => "0000000000000000", 30003 => "0000000000000000", 30004 => "0000000000000000", 30005 => "0000000000000000", 30006 => "0000000000000000", 30007 => "0000000000000000", 30008 => "0000000000000000", 30009 => "0000000000000000", 30010 => "0000000000000000", 30011 => "0000000000000000", 30012 => "0000000000000000", 30013 => "0000000000000000", 30014 => "0000000000000000", 30015 => "0000000000000000", 30016 => "0000000000000000", 30017 => "0000000000000000", 30018 => "0000000000000000", 30019 => "0000000000000000", 30020 => "0000000000000000", 30021 => "0000000000000000", 30022 => "0000000000000000", 30023 => "0000000000000000", 30024 => "0000000000000000", 30025 => "0000000000000000", 30026 => "0000000000000000", 30027 => "0000000000000000", 30028 => "0000000000000000", 30029 => "0000000000000000", 30030 => "0000000000000000", 30031 => "0000000000000000", 30032 => "0000000000000000", 30033 => "0000000000000000", 30034 => "0000000000000000", 30035 => "0000000000000000", 30036 => "0000000000000000", 30037 => "0000000000000000", 30038 => "0000000000000000", 30039 => "0000000000000000", 30040 => "0000000000000000", 30041 => "0000000000000000", 30042 => "0000000000000000", 30043 => "0000000000000000", 30044 => "0000000000000000", 30045 => "0000000000000000", 30046 => "0000000000000000", 30047 => "0000000000000000", 30048 => "0000000000000000", 30049 => "0000000000000000", 30050 => "0000000000000000", 30051 => "0000000000000000", 30052 => "0000000000000000", 30053 => "0000000000000000", 30054 => "0000000000000000", 30055 => "0000000000000000", 30056 => "0000000000000000", 30057 => "0000000000000000", 30058 => "0000000000000000", 30059 => "0000000000000000", 30060 => "0000000000000000", 30061 => "0000000000000000", 30062 => "0000000000000000", 30063 => "0000000000000000", 30064 => "0000000000000000", 30065 => "0000000000000000", 30066 => "0000000000000000", 30067 => "0000000000000000", 30068 => "0000000000000000", 30069 => "0000000000000000", 30070 => "0000000000000000", 30071 => "0000000000000000", 30072 => "0000000000000000", 30073 => "0000000000000000", 30074 => "0000000000000000", 30075 => "0000000000000000", 30076 => "0000000000000000", 30077 => "0000000000000000", 30078 => "0000000000000000", 30079 => "0000000000000000", 30080 => "0000000000000000", 30081 => "0000000000000000", 30082 => "0000000000000000", 30083 => "0000000000000000", 30084 => "0000000000000000", 30085 => "0000000000000000", 30086 => "0000000000000000", 30087 => "0000000000000000", 30088 => "0000000000000000", 30089 => "0000000000000000", 30090 => "0000000000000000", 30091 => "0000000000000000", 30092 => "0000000000000000", 30093 => "0000000000000000", 30094 => "0000000000000000", 30095 => "0000000000000000", 30096 => "0000000000000000", 30097 => "0000000000000000", 30098 => "0000000000000000", 30099 => "0000000000000000", 30100 => "0000000000000000", 30101 => "0000000000000000", 30102 => "0000000000000000", 30103 => "0000000000000000", 30104 => "0000000000000000", 30105 => "0000000000000000", 30106 => "0000000000000000", 30107 => "0000000000000000", 30108 => "0000000000000000", 30109 => "0000000000000000", 30110 => "0000000000000000", 30111 => "0000000000000000", 30112 => "0000000000000000", 30113 => "0000000000000000", 30114 => "0000000000000000", 30115 => "0000000000000000", 30116 => "0000000000000000", 30117 => "0000000000000000", 30118 => "0000000000000000", 30119 => "0000000000000000", 30120 => "0000000000000000", 30121 => "0000000000000000", 30122 => "0000000000000000", 30123 => "0000000000000000", 30124 => "0000000000000000", 30125 => "0000000000000000", 30126 => "0000000000000000", 30127 => "0000000000000000", 30128 => "0000000000000000", 30129 => "0000000000000000", 30130 => "0000000000000000", 30131 => "0000000000000000", 30132 => "0000000000000000", 30133 => "0000000000000000", 30134 => "0000000000000000", 30135 => "0000000000000000", 30136 => "0000000000000000", 30137 => "0000000000000000", 30138 => "0000000000000000", 30139 => "0000000000000000", 30140 => "0000000000000000", 30141 => "0000000000000000", 30142 => "0000000000000000", 30143 => "0000000000000000", 30144 => "0000000000000000", 30145 => "0000000000000000", 30146 => "0000000000000000", 30147 => "0000000000000000", 30148 => "0000000000000000", 30149 => "0000000000000000", 30150 => "0000000000000000", 30151 => "0000000000000000", 30152 => "0000000000000000", 30153 => "0000000000000000", 30154 => "0000000000000000", 30155 => "0000000000000000", 30156 => "0000000000000000", 30157 => "0000000000000000", 30158 => "0000000000000000", 30159 => "0000000000000000", 30160 => "0000000000000000", 30161 => "0000000000000000", 30162 => "0000000000000000", 30163 => "0000000000000000", 30164 => "0000000000000000", 30165 => "0000000000000000", 30166 => "0000000000000000", 30167 => "0000000000000000", 30168 => "0000000000000000", 30169 => "0000000000000000", 30170 => "0000000000000000", 30171 => "0000000000000000", 30172 => "0000000000000000", 30173 => "0000000000000000", 30174 => "0000000000000000", 30175 => "0000000000000000", 30176 => "0000000000000000", 30177 => "0000000000000000", 30178 => "0000000000000000", 30179 => "0000000000000000", 30180 => "0000000000000000", 30181 => "0000000000000000", 30182 => "0000000000000000", 30183 => "0000000000000000", 30184 => "0000000000000000", 30185 => "0000000000000000", 30186 => "0000000000000000", 30187 => "0000000000000000", 30188 => "0000000000000000", 30189 => "0000000000000000", 30190 => "0000000000000000", 30191 => "0000000000000000", 30192 => "0000000000000000", 30193 => "0000000000000000", 30194 => "0000000000000000", 30195 => "0000000000000000", 30196 => "0000000000000000", 30197 => "0000000000000000", 30198 => "0000000000000000", 30199 => "0000000000000000", 30200 => "0000000000000000", 30201 => "0000000000000000", 30202 => "0000000000000000", 30203 => "0000000000000000", 30204 => "0000000000000000", 30205 => "0000000000000000", 30206 => "0000000000000000", 30207 => "0000000000000000", 30208 => "0000000000000000", 30209 => "0000000000000000", 30210 => "0000000000000000", 30211 => "0000000000000000", 30212 => "0000000000000000", 30213 => "0000000000000000", 30214 => "0000000000000000", 30215 => "0000000000000000", 30216 => "0000000000000000", 30217 => "0000000000000000", 30218 => "0000000000000000", 30219 => "0000000000000000", 30220 => "0000000000000000", 30221 => "0000000000000000", 30222 => "0000000000000000", 30223 => "0000000000000000", 30224 => "0000000000000000", 30225 => "0000000000000000", 30226 => "0000000000000000", 30227 => "0000000000000000", 30228 => "0000000000000000", 30229 => "0000000000000000", 30230 => "0000000000000000", 30231 => "0000000000000000", 30232 => "0000000000000000", 30233 => "0000000000000000", 30234 => "0000000000000000", 30235 => "0000000000000000", 30236 => "0000000000000000", 30237 => "0000000000000000", 30238 => "0000000000000000", 30239 => "0000000000000000", 30240 => "0000000000000000", 30241 => "0000000000000000", 30242 => "0000000000000000", 30243 => "0000000000000000", 30244 => "0000000000000000", 30245 => "0000000000000000", 30246 => "0000000000000000", 30247 => "0000000000000000", 30248 => "0000000000000000", 30249 => "0000000000000000", 30250 => "0000000000000000", 30251 => "0000000000000000", 30252 => "0000000000000000", 30253 => "0000000000000000", 30254 => "0000000000000000", 30255 => "0000000000000000", 30256 => "0000000000000000", 30257 => "0000000000000000", 30258 => "0000000000000000", 30259 => "0000000000000000", 30260 => "0000000000000000", 30261 => "0000000000000000", 30262 => "0000000000000000", 30263 => "0000000000000000", 30264 => "0000000000000000", 30265 => "0000000000000000", 30266 => "0000000000000000", 30267 => "0000000000000000", 30268 => "0000000000000000", 30269 => "0000000000000000", 30270 => "0000000000000000", 30271 => "0000000000000000", 30272 => "0000000000000000", 30273 => "0000000000000000", 30274 => "0000000000000000", 30275 => "0000000000000000", 30276 => "0000000000000000", 30277 => "0000000000000000", 30278 => "0000000000000000", 30279 => "0000000000000000", 30280 => "0000000000000000", 30281 => "0000000000000000", 30282 => "0000000000000000", 30283 => "0000000000000000", 30284 => "0000000000000000", 30285 => "0000000000000000", 30286 => "0000000000000000", 30287 => "0000000000000000", 30288 => "0000000000000000", 30289 => "0000000000000000", 30290 => "0000000000000000", 30291 => "0000000000000000", 30292 => "0000000000000000", 30293 => "0000000000000000", 30294 => "0000000000000000", 30295 => "0000000000000000", 30296 => "0000000000000000", 30297 => "0000000000000000", 30298 => "0000000000000000", 30299 => "0000000000000000", 30300 => "0000000000000000", 30301 => "0000000000000000", 30302 => "0000000000000000", 30303 => "0000000000000000", 30304 => "0000000000000000", 30305 => "0000000000000000", 30306 => "0000000000000000", 30307 => "0000000000000000", 30308 => "0000000000000000", 30309 => "0000000000000000", 30310 => "0000000000000000", 30311 => "0000000000000000", 30312 => "0000000000000000", 30313 => "0000000000000000", 30314 => "0000000000000000", 30315 => "0000000000000000", 30316 => "0000000000000000", 30317 => "0000000000000000", 30318 => "0000000000000000", 30319 => "0000000000000000", 30320 => "0000000000000000", 30321 => "0000000000000000", 30322 => "0000000000000000", 30323 => "0000000000000000", 30324 => "0000000000000000", 30325 => "0000000000000000", 30326 => "0000000000000000", 30327 => "0000000000000000", 30328 => "0000000000000000", 30329 => "0000000000000000", 30330 => "0000000000000000", 30331 => "0000000000000000", 30332 => "0000000000000000", 30333 => "0000000000000000", 30334 => "0000000000000000", 30335 => "0000000000000000", 30336 => "0000000000000000", 30337 => "0000000000000000", 30338 => "0000000000000000", 30339 => "0000000000000000", 30340 => "0000000000000000", 30341 => "0000000000000000", 30342 => "0000000000000000", 30343 => "0000000000000000", 30344 => "0000000000000000", 30345 => "0000000000000000", 30346 => "0000000000000000", 30347 => "0000000000000000", 30348 => "0000000000000000", 30349 => "0000000000000000", 30350 => "0000000000000000", 30351 => "0000000000000000", 30352 => "0000000000000000", 30353 => "0000000000000000", 30354 => "0000000000000000", 30355 => "0000000000000000", 30356 => "0000000000000000", 30357 => "0000000000000000", 30358 => "0000000000000000", 30359 => "0000000000000000", 30360 => "0000000000000000", 30361 => "0000000000000000", 30362 => "0000000000000000", 30363 => "0000000000000000", 30364 => "0000000000000000", 30365 => "0000000000000000", 30366 => "0000000000000000", 30367 => "0000000000000000", 30368 => "0000000000000000", 30369 => "0000000000000000", 30370 => "0000000000000000", 30371 => "0000000000000000", 30372 => "0000000000000000", 30373 => "0000000000000000", 30374 => "0000000000000000", 30375 => "0000000000000000", 30376 => "0000000000000000", 30377 => "0000000000000000", 30378 => "0000000000000000", 30379 => "0000000000000000", 30380 => "0000000000000000", 30381 => "0000000000000000", 30382 => "0000000000000000", 30383 => "0000000000000000", 30384 => "0000000000000000", 30385 => "0000000000000000", 30386 => "0000000000000000", 30387 => "0000000000000000", 30388 => "0000000000000000", 30389 => "0000000000000000", 30390 => "0000000000000000", 30391 => "0000000000000000", 30392 => "0000000000000000", 30393 => "0000000000000000", 30394 => "0000000000000000", 30395 => "0000000000000000", 30396 => "0000000000000000", 30397 => "0000000000000000", 30398 => "0000000000000000", 30399 => "0000000000000000", 30400 => "0000000000000000", 30401 => "0000000000000000", 30402 => "0000000000000000", 30403 => "0000000000000000", 30404 => "0000000000000000", 30405 => "0000000000000000", 30406 => "0000000000000000", 30407 => "0000000000000000", 30408 => "0000000000000000", 30409 => "0000000000000000", 30410 => "0000000000000000", 30411 => "0000000000000000", 30412 => "0000000000000000", 30413 => "0000000000000000", 30414 => "0000000000000000", 30415 => "0000000000000000", 30416 => "0000000000000000", 30417 => "0000000000000000", 30418 => "0000000000000000", 30419 => "0000000000000000", 30420 => "0000000000000000", 30421 => "0000000000000000", 30422 => "0000000000000000", 30423 => "0000000000000000", 30424 => "0000000000000000", 30425 => "0000000000000000", 30426 => "0000000000000000", 30427 => "0000000000000000", 30428 => "0000000000000000", 30429 => "0000000000000000", 30430 => "0000000000000000", 30431 => "0000000000000000", 30432 => "0000000000000000", 30433 => "0000000000000000", 30434 => "0000000000000000", 30435 => "0000000000000000", 30436 => "0000000000000000", 30437 => "0000000000000000", 30438 => "0000000000000000", 30439 => "0000000000000000", 30440 => "0000000000000000", 30441 => "0000000000000000", 30442 => "0000000000000000", 30443 => "0000000000000000", 30444 => "0000000000000000", 30445 => "0000000000000000", 30446 => "0000000000000000", 30447 => "0000000000000000", 30448 => "0000000000000000", 30449 => "0000000000000000", 30450 => "0000000000000000", 30451 => "0000000000000000", 30452 => "0000000000000000", 30453 => "0000000000000000", 30454 => "0000000000000000", 30455 => "0000000000000000", 30456 => "0000000000000000", 30457 => "0000000000000000", 30458 => "0000000000000000", 30459 => "0000000000000000", 30460 => "0000000000000000", 30461 => "0000000000000000", 30462 => "0000000000000000", 30463 => "0000000000000000", 30464 => "0000000000000000", 30465 => "0000000000000000", 30466 => "0000000000000000", 30467 => "0000000000000000", 30468 => "0000000000000000", 30469 => "0000000000000000", 30470 => "0000000000000000", 30471 => "0000000000000000", 30472 => "0000000000000000", 30473 => "0000000000000000", 30474 => "0000000000000000", 30475 => "0000000000000000", 30476 => "0000000000000000", 30477 => "0000000000000000", 30478 => "0000000000000000", 30479 => "0000000000000000", 30480 => "0000000000000000", 30481 => "0000000000000000", 30482 => "0000000000000000", 30483 => "0000000000000000", 30484 => "0000000000000000", 30485 => "0000000000000000", 30486 => "0000000000000000", 30487 => "0000000000000000", 30488 => "0000000000000000", 30489 => "0000000000000000", 30490 => "0000000000000000", 30491 => "0000000000000000", 30492 => "0000000000000000", 30493 => "0000000000000000", 30494 => "0000000000000000", 30495 => "0000000000000000", 30496 => "0000000000000000", 30497 => "0000000000000000", 30498 => "0000000000000000", 30499 => "0000000000000000", 30500 => "0000000000000000", 30501 => "0000000000000000", 30502 => "0000000000000000", 30503 => "0000000000000000", 30504 => "0000000000000000", 30505 => "0000000000000000", 30506 => "0000000000000000", 30507 => "0000000000000000", 30508 => "0000000000000000", 30509 => "0000000000000000", 30510 => "0000000000000000", 30511 => "0000000000000000", 30512 => "0000000000000000", 30513 => "0000000000000000", 30514 => "0000000000000000", 30515 => "0000000000000000", 30516 => "0000000000000000", 30517 => "0000000000000000", 30518 => "0000000000000000", 30519 => "0000000000000000", 30520 => "0000000000000000", 30521 => "0000000000000000", 30522 => "0000000000000000", 30523 => "0000000000000000", 30524 => "0000000000000000", 30525 => "0000000000000000", 30526 => "0000000000000000", 30527 => "0000000000000000", 30528 => "0000000000000000", 30529 => "0000000000000000", 30530 => "0000000000000000", 30531 => "0000000000000000", 30532 => "0000000000000000", 30533 => "0000000000000000", 30534 => "0000000000000000", 30535 => "0000000000000000", 30536 => "0000000000000000", 30537 => "0000000000000000", 30538 => "0000000000000000", 30539 => "0000000000000000", 30540 => "0000000000000000", 30541 => "0000000000000000", 30542 => "0000000000000000", 30543 => "0000000000000000", 30544 => "0000000000000000", 30545 => "0000000000000000", 30546 => "0000000000000000", 30547 => "0000000000000000", 30548 => "0000000000000000", 30549 => "0000000000000000", 30550 => "0000000000000000", 30551 => "0000000000000000", 30552 => "0000000000000000", 30553 => "0000000000000000", 30554 => "0000000000000000", 30555 => "0000000000000000", 30556 => "0000000000000000", 30557 => "0000000000000000", 30558 => "0000000000000000", 30559 => "0000000000000000", 30560 => "0000000000000000", 30561 => "0000000000000000", 30562 => "0000000000000000", 30563 => "0000000000000000", 30564 => "0000000000000000", 30565 => "0000000000000000", 30566 => "0000000000000000", 30567 => "0000000000000000", 30568 => "0000000000000000", 30569 => "0000000000000000", 30570 => "0000000000000000", 30571 => "0000000000000000", 30572 => "0000000000000000", 30573 => "0000000000000000", 30574 => "0000000000000000", 30575 => "0000000000000000", 30576 => "0000000000000000", 30577 => "0000000000000000", 30578 => "0000000000000000", 30579 => "0000000000000000", 30580 => "0000000000000000", 30581 => "0000000000000000", 30582 => "0000000000000000", 30583 => "0000000000000000", 30584 => "0000000000000000", 30585 => "0000000000000000", 30586 => "0000000000000000", 30587 => "0000000000000000", 30588 => "0000000000000000", 30589 => "0000000000000000", 30590 => "0000000000000000", 30591 => "0000000000000000", 30592 => "0000000000000000", 30593 => "0000000000000000", 30594 => "0000000000000000", 30595 => "0000000000000000", 30596 => "0000000000000000", 30597 => "0000000000000000", 30598 => "0000000000000000", 30599 => "0000000000000000", 30600 => "0000000000000000", 30601 => "0000000000000000", 30602 => "0000000000000000", 30603 => "0000000000000000", 30604 => "0000000000000000", 30605 => "0000000000000000", 30606 => "0000000000000000", 30607 => "0000000000000000", 30608 => "0000000000000000", 30609 => "0000000000000000", 30610 => "0000000000000000", 30611 => "0000000000000000", 30612 => "0000000000000000", 30613 => "0000000000000000", 30614 => "0000000000000000", 30615 => "0000000000000000", 30616 => "0000000000000000", 30617 => "0000000000000000", 30618 => "0000000000000000", 30619 => "0000000000000000", 30620 => "0000000000000000", 30621 => "0000000000000000", 30622 => "0000000000000000", 30623 => "0000000000000000", 30624 => "0000000000000000", 30625 => "0000000000000000", 30626 => "0000000000000000", 30627 => "0000000000000000", 30628 => "0000000000000000", 30629 => "0000000000000000", 30630 => "0000000000000000", 30631 => "0000000000000000", 30632 => "0000000000000000", 30633 => "0000000000000000", 30634 => "0000000000000000", 30635 => "0000000000000000", 30636 => "0000000000000000", 30637 => "0000000000000000", 30638 => "0000000000000000", 30639 => "0000000000000000", 30640 => "0000000000000000", 30641 => "0000000000000000", 30642 => "0000000000000000", 30643 => "0000000000000000", 30644 => "0000000000000000", 30645 => "0000000000000000", 30646 => "0000000000000000", 30647 => "0000000000000000", 30648 => "0000000000000000", 30649 => "0000000000000000", 30650 => "0000000000000000", 30651 => "0000000000000000", 30652 => "0000000000000000", 30653 => "0000000000000000", 30654 => "0000000000000000", 30655 => "0000000000000000", 30656 => "0000000000000000", 30657 => "0000000000000000", 30658 => "0000000000000000", 30659 => "0000000000000000", 30660 => "0000000000000000", 30661 => "0000000000000000", 30662 => "0000000000000000", 30663 => "0000000000000000", 30664 => "0000000000000000", 30665 => "0000000000000000", 30666 => "0000000000000000", 30667 => "0000000000000000", 30668 => "0000000000000000", 30669 => "0000000000000000", 30670 => "0000000000000000", 30671 => "0000000000000000", 30672 => "0000000000000000", 30673 => "0000000000000000", 30674 => "0000000000000000", 30675 => "0000000000000000", 30676 => "0000000000000000", 30677 => "0000000000000000", 30678 => "0000000000000000", 30679 => "0000000000000000", 30680 => "0000000000000000", 30681 => "0000000000000000", 30682 => "0000000000000000", 30683 => "0000000000000000", 30684 => "0000000000000000", 30685 => "0000000000000000", 30686 => "0000000000000000", 30687 => "0000000000000000", 30688 => "0000000000000000", 30689 => "0000000000000000", 30690 => "0000000000000000", 30691 => "0000000000000000", 30692 => "0000000000000000", 30693 => "0000000000000000", 30694 => "0000000000000000", 30695 => "0000000000000000", 30696 => "0000000000000000", 30697 => "0000000000000000", 30698 => "0000000000000000", 30699 => "0000000000000000", 30700 => "0000000000000000", 30701 => "0000000000000000", 30702 => "0000000000000000", 30703 => "0000000000000000", 30704 => "0000000000000000", 30705 => "0000000000000000", 30706 => "0000000000000000", 30707 => "0000000000000000", 30708 => "0000000000000000", 30709 => "0000000000000000", 30710 => "0000000000000000", 30711 => "0000000000000000", 30712 => "0000000000000000", 30713 => "0000000000000000", 30714 => "0000000000000000", 30715 => "0000000000000000", 30716 => "0000000000000000", 30717 => "0000000000000000", 30718 => "0000000000000000", 30719 => "0000000000000000", 30720 => "0000000000000000", 30721 => "0000000000000000", 30722 => "0000000000000000", 30723 => "0000000000000000", 30724 => "0000000000000000", 30725 => "0000000000000000", 30726 => "0000000000000000", 30727 => "0000000000000000", 30728 => "0000000000000000", 30729 => "0000000000000000", 30730 => "0000000000000000", 30731 => "0000000000000000", 30732 => "0000000000000000", 30733 => "0000000000000000", 30734 => "0000000000000000", 30735 => "0000000000000000", 30736 => "0000000000000000", 30737 => "0000000000000000", 30738 => "0000000000000000", 30739 => "0000000000000000", 30740 => "0000000000000000", 30741 => "0000000000000000", 30742 => "0000000000000000", 30743 => "0000000000000000", 30744 => "0000000000000000", 30745 => "0000000000000000", 30746 => "0000000000000000", 30747 => "0000000000000000", 30748 => "0000000000000000", 30749 => "0000000000000000", 30750 => "0000000000000000", 30751 => "0000000000000000", 30752 => "0000000000000000", 30753 => "0000000000000000", 30754 => "0000000000000000", 30755 => "0000000000000000", 30756 => "0000000000000000", 30757 => "0000000000000000", 30758 => "0000000000000000", 30759 => "0000000000000000", 30760 => "0000000000000000", 30761 => "0000000000000000", 30762 => "0000000000000000", 30763 => "0000000000000000", 30764 => "0000000000000000", 30765 => "0000000000000000", 30766 => "0000000000000000", 30767 => "0000000000000000", 30768 => "0000000000000000", 30769 => "0000000000000000", 30770 => "0000000000000000", 30771 => "0000000000000000", 30772 => "0000000000000000", 30773 => "0000000000000000", 30774 => "0000000000000000", 30775 => "0000000000000000", 30776 => "0000000000000000", 30777 => "0000000000000000", 30778 => "0000000000000000", 30779 => "0000000000000000", 30780 => "0000000000000000", 30781 => "0000000000000000", 30782 => "0000000000000000", 30783 => "0000000000000000", 30784 => "0000000000000000", 30785 => "0000000000000000", 30786 => "0000000000000000", 30787 => "0000000000000000", 30788 => "0000000000000000", 30789 => "0000000000000000", 30790 => "0000000000000000", 30791 => "0000000000000000", 30792 => "0000000000000000", 30793 => "0000000000000000", 30794 => "0000000000000000", 30795 => "0000000000000000", 30796 => "0000000000000000", 30797 => "0000000000000000", 30798 => "0000000000000000", 30799 => "0000000000000000", 30800 => "0000000000000000", 30801 => "0000000000000000", 30802 => "0000000000000000", 30803 => "0000000000000000", 30804 => "0000000000000000", 30805 => "0000000000000000", 30806 => "0000000000000000", 30807 => "0000000000000000", 30808 => "0000000000000000", 30809 => "0000000000000000", 30810 => "0000000000000000", 30811 => "0000000000000000", 30812 => "0000000000000000", 30813 => "0000000000000000", 30814 => "0000000000000000", 30815 => "0000000000000000", 30816 => "0000000000000000", 30817 => "0000000000000000", 30818 => "0000000000000000", 30819 => "0000000000000000", 30820 => "0000000000000000", 30821 => "0000000000000000", 30822 => "0000000000000000", 30823 => "0000000000000000", 30824 => "0000000000000000", 30825 => "0000000000000000", 30826 => "0000000000000000", 30827 => "0000000000000000", 30828 => "0000000000000000", 30829 => "0000000000000000", 30830 => "0000000000000000", 30831 => "0000000000000000", 30832 => "0000000000000000", 30833 => "0000000000000000", 30834 => "0000000000000000", 30835 => "0000000000000000", 30836 => "0000000000000000", 30837 => "0000000000000000", 30838 => "0000000000000000", 30839 => "0000000000000000", 30840 => "0000000000000000", 30841 => "0000000000000000", 30842 => "0000000000000000", 30843 => "0000000000000000", 30844 => "0000000000000000", 30845 => "0000000000000000", 30846 => "0000000000000000", 30847 => "0000000000000000", 30848 => "0000000000000000", 30849 => "0000000000000000", 30850 => "0000000000000000", 30851 => "0000000000000000", 30852 => "0000000000000000", 30853 => "0000000000000000", 30854 => "0000000000000000", 30855 => "0000000000000000", 30856 => "0000000000000000", 30857 => "0000000000000000", 30858 => "0000000000000000", 30859 => "0000000000000000", 30860 => "0000000000000000", 30861 => "0000000000000000", 30862 => "0000000000000000", 30863 => "0000000000000000", 30864 => "0000000000000000", 30865 => "0000000000000000", 30866 => "0000000000000000", 30867 => "0000000000000000", 30868 => "0000000000000000", 30869 => "0000000000000000", 30870 => "0000000000000000", 30871 => "0000000000000000", 30872 => "0000000000000000", 30873 => "0000000000000000", 30874 => "0000000000000000", 30875 => "0000000000000000", 30876 => "0000000000000000", 30877 => "0000000000000000", 30878 => "0000000000000000", 30879 => "0000000000000000", 30880 => "0000000000000000", 30881 => "0000000000000000", 30882 => "0000000000000000", 30883 => "0000000000000000", 30884 => "0000000000000000", 30885 => "0000000000000000", 30886 => "0000000000000000", 30887 => "0000000000000000", 30888 => "0000000000000000", 30889 => "0000000000000000", 30890 => "0000000000000000", 30891 => "0000000000000000", 30892 => "0000000000000000", 30893 => "0000000000000000", 30894 => "0000000000000000", 30895 => "0000000000000000", 30896 => "0000000000000000", 30897 => "0000000000000000", 30898 => "0000000000000000", 30899 => "0000000000000000", 30900 => "0000000000000000", 30901 => "0000000000000000", 30902 => "0000000000000000", 30903 => "0000000000000000", 30904 => "0000000000000000", 30905 => "0000000000000000", 30906 => "0000000000000000", 30907 => "0000000000000000", 30908 => "0000000000000000", 30909 => "0000000000000000", 30910 => "0000000000000000", 30911 => "0000000000000000", 30912 => "0000000000000000", 30913 => "0000000000000000", 30914 => "0000000000000000", 30915 => "0000000000000000", 30916 => "0000000000000000", 30917 => "0000000000000000", 30918 => "0000000000000000", 30919 => "0000000000000000", 30920 => "0000000000000000", 30921 => "0000000000000000", 30922 => "0000000000000000", 30923 => "0000000000000000", 30924 => "0000000000000000", 30925 => "0000000000000000", 30926 => "0000000000000000", 30927 => "0000000000000000", 30928 => "0000000000000000", 30929 => "0000000000000000", 30930 => "0000000000000000", 30931 => "0000000000000000", 30932 => "0000000000000000", 30933 => "0000000000000000", 30934 => "0000000000000000", 30935 => "0000000000000000", 30936 => "0000000000000000", 30937 => "0000000000000000", 30938 => "0000000000000000", 30939 => "0000000000000000", 30940 => "0000000000000000", 30941 => "0000000000000000", 30942 => "0000000000000000", 30943 => "0000000000000000", 30944 => "0000000000000000", 30945 => "0000000000000000", 30946 => "0000000000000000", 30947 => "0000000000000000", 30948 => "0000000000000000", 30949 => "0000000000000000", 30950 => "0000000000000000", 30951 => "0000000000000000", 30952 => "0000000000000000", 30953 => "0000000000000000", 30954 => "0000000000000000", 30955 => "0000000000000000", 30956 => "0000000000000000", 30957 => "0000000000000000", 30958 => "0000000000000000", 30959 => "0000000000000000", 30960 => "0000000000000000", 30961 => "0000000000000000", 30962 => "0000000000000000", 30963 => "0000000000000000", 30964 => "0000000000000000", 30965 => "0000000000000000", 30966 => "0000000000000000", 30967 => "0000000000000000", 30968 => "0000000000000000", 30969 => "0000000000000000", 30970 => "0000000000000000", 30971 => "0000000000000000", 30972 => "0000000000000000", 30973 => "0000000000000000", 30974 => "0000000000000000", 30975 => "0000000000000000", 30976 => "0000000000000000", 30977 => "0000000000000000", 30978 => "0000000000000000", 30979 => "0000000000000000", 30980 => "0000000000000000", 30981 => "0000000000000000", 30982 => "0000000000000000", 30983 => "0000000000000000", 30984 => "0000000000000000", 30985 => "0000000000000000", 30986 => "0000000000000000", 30987 => "0000000000000000", 30988 => "0000000000000000", 30989 => "0000000000000000", 30990 => "0000000000000000", 30991 => "0000000000000000", 30992 => "0000000000000000", 30993 => "0000000000000000", 30994 => "0000000000000000", 30995 => "0000000000000000", 30996 => "0000000000000000", 30997 => "0000000000000000", 30998 => "0000000000000000", 30999 => "0000000000000000", 31000 => "0000000000000000", 31001 => "0000000000000000", 31002 => "0000000000000000", 31003 => "0000000000000000", 31004 => "0000000000000000", 31005 => "0000000000000000", 31006 => "0000000000000000", 31007 => "0000000000000000", 31008 => "0000000000000000", 31009 => "0000000000000000", 31010 => "0000000000000000", 31011 => "0000000000000000", 31012 => "0000000000000000", 31013 => "0000000000000000", 31014 => "0000000000000000", 31015 => "0000000000000000", 31016 => "0000000000000000", 31017 => "0000000000000000", 31018 => "0000000000000000", 31019 => "0000000000000000", 31020 => "0000000000000000", 31021 => "0000000000000000", 31022 => "0000000000000000", 31023 => "0000000000000000", 31024 => "0000000000000000", 31025 => "0000000000000000", 31026 => "0000000000000000", 31027 => "0000000000000000", 31028 => "0000000000000000", 31029 => "0000000000000000", 31030 => "0000000000000000", 31031 => "0000000000000000", 31032 => "0000000000000000", 31033 => "0000000000000000", 31034 => "0000000000000000", 31035 => "0000000000000000", 31036 => "0000000000000000", 31037 => "0000000000000000", 31038 => "0000000000000000", 31039 => "0000000000000000", 31040 => "0000000000000000", 31041 => "0000000000000000", 31042 => "0000000000000000", 31043 => "0000000000000000", 31044 => "0000000000000000", 31045 => "0000000000000000", 31046 => "0000000000000000", 31047 => "0000000000000000", 31048 => "0000000000000000", 31049 => "0000000000000000", 31050 => "0000000000000000", 31051 => "0000000000000000", 31052 => "0000000000000000", 31053 => "0000000000000000", 31054 => "0000000000000000", 31055 => "0000000000000000", 31056 => "0000000000000000", 31057 => "0000000000000000", 31058 => "0000000000000000", 31059 => "0000000000000000", 31060 => "0000000000000000", 31061 => "0000000000000000", 31062 => "0000000000000000", 31063 => "0000000000000000", 31064 => "0000000000000000", 31065 => "0000000000000000", 31066 => "0000000000000000", 31067 => "0000000000000000", 31068 => "0000000000000000", 31069 => "0000000000000000", 31070 => "0000000000000000", 31071 => "0000000000000000", 31072 => "0000000000000000", 31073 => "0000000000000000", 31074 => "0000000000000000", 31075 => "0000000000000000", 31076 => "0000000000000000", 31077 => "0000000000000000", 31078 => "0000000000000000", 31079 => "0000000000000000", 31080 => "0000000000000000", 31081 => "0000000000000000", 31082 => "0000000000000000", 31083 => "0000000000000000", 31084 => "0000000000000000", 31085 => "0000000000000000", 31086 => "0000000000000000", 31087 => "0000000000000000", 31088 => "0000000000000000", 31089 => "0000000000000000", 31090 => "0000000000000000", 31091 => "0000000000000000", 31092 => "0000000000000000", 31093 => "0000000000000000", 31094 => "0000000000000000", 31095 => "0000000000000000", 31096 => "0000000000000000", 31097 => "0000000000000000", 31098 => "0000000000000000", 31099 => "0000000000000000", 31100 => "0000000000000000", 31101 => "0000000000000000", 31102 => "0000000000000000", 31103 => "0000000000000000", 31104 => "0000000000000000", 31105 => "0000000000000000", 31106 => "0000000000000000", 31107 => "0000000000000000", 31108 => "0000000000000000", 31109 => "0000000000000000", 31110 => "0000000000000000", 31111 => "0000000000000000", 31112 => "0000000000000000", 31113 => "0000000000000000", 31114 => "0000000000000000", 31115 => "0000000000000000", 31116 => "0000000000000000", 31117 => "0000000000000000", 31118 => "0000000000000000", 31119 => "0000000000000000", 31120 => "0000000000000000", 31121 => "0000000000000000", 31122 => "0000000000000000", 31123 => "0000000000000000", 31124 => "0000000000000000", 31125 => "0000000000000000", 31126 => "0000000000000000", 31127 => "0000000000000000", 31128 => "0000000000000000", 31129 => "0000000000000000", 31130 => "0000000000000000", 31131 => "0000000000000000", 31132 => "0000000000000000", 31133 => "0000000000000000", 31134 => "0000000000000000", 31135 => "0000000000000000", 31136 => "0000000000000000", 31137 => "0000000000000000", 31138 => "0000000000000000", 31139 => "0000000000000000", 31140 => "0000000000000000", 31141 => "0000000000000000", 31142 => "0000000000000000", 31143 => "0000000000000000", 31144 => "0000000000000000", 31145 => "0000000000000000", 31146 => "0000000000000000", 31147 => "0000000000000000", 31148 => "0000000000000000", 31149 => "0000000000000000", 31150 => "0000000000000000", 31151 => "0000000000000000", 31152 => "0000000000000000", 31153 => "0000000000000000", 31154 => "0000000000000000", 31155 => "0000000000000000", 31156 => "0000000000000000", 31157 => "0000000000000000", 31158 => "0000000000000000", 31159 => "0000000000000000", 31160 => "0000000000000000", 31161 => "0000000000000000", 31162 => "0000000000000000", 31163 => "0000000000000000", 31164 => "0000000000000000", 31165 => "0000000000000000", 31166 => "0000000000000000", 31167 => "0000000000000000", 31168 => "0000000000000000", 31169 => "0000000000000000", 31170 => "0000000000000000", 31171 => "0000000000000000", 31172 => "0000000000000000", 31173 => "0000000000000000", 31174 => "0000000000000000", 31175 => "0000000000000000", 31176 => "0000000000000000", 31177 => "0000000000000000", 31178 => "0000000000000000", 31179 => "0000000000000000", 31180 => "0000000000000000", 31181 => "0000000000000000", 31182 => "0000000000000000", 31183 => "0000000000000000", 31184 => "0000000000000000", 31185 => "0000000000000000", 31186 => "0000000000000000", 31187 => "0000000000000000", 31188 => "0000000000000000", 31189 => "0000000000000000", 31190 => "0000000000000000", 31191 => "0000000000000000", 31192 => "0000000000000000", 31193 => "0000000000000000", 31194 => "0000000000000000", 31195 => "0000000000000000", 31196 => "0000000000000000", 31197 => "0000000000000000", 31198 => "0000000000000000", 31199 => "0000000000000000", 31200 => "0000000000000000", 31201 => "0000000000000000", 31202 => "0000000000000000", 31203 => "0000000000000000", 31204 => "0000000000000000", 31205 => "0000000000000000", 31206 => "0000000000000000", 31207 => "0000000000000000", 31208 => "0000000000000000", 31209 => "0000000000000000", 31210 => "0000000000000000", 31211 => "0000000000000000", 31212 => "0000000000000000", 31213 => "0000000000000000", 31214 => "0000000000000000", 31215 => "0000000000000000", 31216 => "0000000000000000", 31217 => "0000000000000000", 31218 => "0000000000000000", 31219 => "0000000000000000", 31220 => "0000000000000000", 31221 => "0000000000000000", 31222 => "0000000000000000", 31223 => "0000000000000000", 31224 => "0000000000000000", 31225 => "0000000000000000", 31226 => "0000000000000000", 31227 => "0000000000000000", 31228 => "0000000000000000", 31229 => "0000000000000000", 31230 => "0000000000000000", 31231 => "0000000000000000", 31232 => "0000000000000000", 31233 => "0000000000000000", 31234 => "0000000000000000", 31235 => "0000000000000000", 31236 => "0000000000000000", 31237 => "0000000000000000", 31238 => "0000000000000000", 31239 => "0000000000000000", 31240 => "0000000000000000", 31241 => "0000000000000000", 31242 => "0000000000000000", 31243 => "0000000000000000", 31244 => "0000000000000000", 31245 => "0000000000000000", 31246 => "0000000000000000", 31247 => "0000000000000000", 31248 => "0000000000000000", 31249 => "0000000000000000", 31250 => "0000000000000000", 31251 => "0000000000000000", 31252 => "0000000000000000", 31253 => "0000000000000000", 31254 => "0000000000000000", 31255 => "0000000000000000", 31256 => "0000000000000000", 31257 => "0000000000000000", 31258 => "0000000000000000", 31259 => "0000000000000000", 31260 => "0000000000000000", 31261 => "0000000000000000", 31262 => "0000000000000000", 31263 => "0000000000000000", 31264 => "0000000000000000", 31265 => "0000000000000000", 31266 => "0000000000000000", 31267 => "0000000000000000", 31268 => "0000000000000000", 31269 => "0000000000000000", 31270 => "0000000000000000", 31271 => "0000000000000000", 31272 => "0000000000000000", 31273 => "0000000000000000", 31274 => "0000000000000000", 31275 => "0000000000000000", 31276 => "0000000000000000", 31277 => "0000000000000000", 31278 => "0000000000000000", 31279 => "0000000000000000", 31280 => "0000000000000000", 31281 => "0000000000000000", 31282 => "0000000000000000", 31283 => "0000000000000000", 31284 => "0000000000000000", 31285 => "0000000000000000", 31286 => "0000000000000000", 31287 => "0000000000000000", 31288 => "0000000000000000", 31289 => "0000000000000000", 31290 => "0000000000000000", 31291 => "0000000000000000", 31292 => "0000000000000000", 31293 => "0000000000000000", 31294 => "0000000000000000", 31295 => "0000000000000000", 31296 => "0000000000000000", 31297 => "0000000000000000", 31298 => "0000000000000000", 31299 => "0000000000000000", 31300 => "0000000000000000", 31301 => "0000000000000000", 31302 => "0000000000000000", 31303 => "0000000000000000", 31304 => "0000000000000000", 31305 => "0000000000000000", 31306 => "0000000000000000", 31307 => "0000000000000000", 31308 => "0000000000000000", 31309 => "0000000000000000", 31310 => "0000000000000000", 31311 => "0000000000000000", 31312 => "0000000000000000", 31313 => "0000000000000000", 31314 => "0000000000000000", 31315 => "0000000000000000", 31316 => "0000000000000000", 31317 => "0000000000000000", 31318 => "0000000000000000", 31319 => "0000000000000000", 31320 => "0000000000000000", 31321 => "0000000000000000", 31322 => "0000000000000000", 31323 => "0000000000000000", 31324 => "0000000000000000", 31325 => "0000000000000000", 31326 => "0000000000000000", 31327 => "0000000000000000", 31328 => "0000000000000000", 31329 => "0000000000000000", 31330 => "0000000000000000", 31331 => "0000000000000000", 31332 => "0000000000000000", 31333 => "0000000000000000", 31334 => "0000000000000000", 31335 => "0000000000000000", 31336 => "0000000000000000", 31337 => "0000000000000000", 31338 => "0000000000000000", 31339 => "0000000000000000", 31340 => "0000000000000000", 31341 => "0000000000000000", 31342 => "0000000000000000", 31343 => "0000000000000000", 31344 => "0000000000000000", 31345 => "0000000000000000", 31346 => "0000000000000000", 31347 => "0000000000000000", 31348 => "0000000000000000", 31349 => "0000000000000000", 31350 => "0000000000000000", 31351 => "0000000000000000", 31352 => "0000000000000000", 31353 => "0000000000000000", 31354 => "0000000000000000", 31355 => "0000000000000000", 31356 => "0000000000000000", 31357 => "0000000000000000", 31358 => "0000000000000000", 31359 => "0000000000000000", 31360 => "0000000000000000", 31361 => "0000000000000000", 31362 => "0000000000000000", 31363 => "0000000000000000", 31364 => "0000000000000000", 31365 => "0000000000000000", 31366 => "0000000000000000", 31367 => "0000000000000000", 31368 => "0000000000000000", 31369 => "0000000000000000", 31370 => "0000000000000000", 31371 => "0000000000000000", 31372 => "0000000000000000", 31373 => "0000000000000000", 31374 => "0000000000000000", 31375 => "0000000000000000", 31376 => "0000000000000000", 31377 => "0000000000000000", 31378 => "0000000000000000", 31379 => "0000000000000000", 31380 => "0000000000000000", 31381 => "0000000000000000", 31382 => "0000000000000000", 31383 => "0000000000000000", 31384 => "0000000000000000", 31385 => "0000000000000000", 31386 => "0000000000000000", 31387 => "0000000000000000", 31388 => "0000000000000000", 31389 => "0000000000000000", 31390 => "0000000000000000", 31391 => "0000000000000000", 31392 => "0000000000000000", 31393 => "0000000000000000", 31394 => "0000000000000000", 31395 => "0000000000000000", 31396 => "0000000000000000", 31397 => "0000000000000000", 31398 => "0000000000000000", 31399 => "0000000000000000", 31400 => "0000000000000000", 31401 => "0000000000000000", 31402 => "0000000000000000", 31403 => "0000000000000000", 31404 => "0000000000000000", 31405 => "0000000000000000", 31406 => "0000000000000000", 31407 => "0000000000000000", 31408 => "0000000000000000", 31409 => "0000000000000000", 31410 => "0000000000000000", 31411 => "0000000000000000", 31412 => "0000000000000000", 31413 => "0000000000000000", 31414 => "0000000000000000", 31415 => "0000000000000000", 31416 => "0000000000000000", 31417 => "0000000000000000", 31418 => "0000000000000000", 31419 => "0000000000000000", 31420 => "0000000000000000", 31421 => "0000000000000000", 31422 => "0000000000000000", 31423 => "0000000000000000", 31424 => "0000000000000000", 31425 => "0000000000000000", 31426 => "0000000000000000", 31427 => "0000000000000000", 31428 => "0000000000000000", 31429 => "0000000000000000", 31430 => "0000000000000000", 31431 => "0000000000000000", 31432 => "0000000000000000", 31433 => "0000000000000000", 31434 => "0000000000000000", 31435 => "0000000000000000", 31436 => "0000000000000000", 31437 => "0000000000000000", 31438 => "0000000000000000", 31439 => "0000000000000000", 31440 => "0000000000000000", 31441 => "0000000000000000", 31442 => "0000000000000000", 31443 => "0000000000000000", 31444 => "0000000000000000", 31445 => "0000000000000000", 31446 => "0000000000000000", 31447 => "0000000000000000", 31448 => "0000000000000000", 31449 => "0000000000000000", 31450 => "0000000000000000", 31451 => "0000000000000000", 31452 => "0000000000000000", 31453 => "0000000000000000", 31454 => "0000000000000000", 31455 => "0000000000000000", 31456 => "0000000000000000", 31457 => "0000000000000000", 31458 => "0000000000000000", 31459 => "0000000000000000", 31460 => "0000000000000000", 31461 => "0000000000000000", 31462 => "0000000000000000", 31463 => "0000000000000000", 31464 => "0000000000000000", 31465 => "0000000000000000", 31466 => "0000000000000000", 31467 => "0000000000000000", 31468 => "0000000000000000", 31469 => "0000000000000000", 31470 => "0000000000000000", 31471 => "0000000000000000", 31472 => "0000000000000000", 31473 => "0000000000000000", 31474 => "0000000000000000", 31475 => "0000000000000000", 31476 => "0000000000000000", 31477 => "0000000000000000", 31478 => "0000000000000000", 31479 => "0000000000000000", 31480 => "0000000000000000", 31481 => "0000000000000000", 31482 => "0000000000000000", 31483 => "0000000000000000", 31484 => "0000000000000000", 31485 => "0000000000000000", 31486 => "0000000000000000", 31487 => "0000000000000000", 31488 => "0000000000000000", 31489 => "0000000000000000", 31490 => "0000000000000000", 31491 => "0000000000000000", 31492 => "0000000000000000", 31493 => "0000000000000000", 31494 => "0000000000000000", 31495 => "0000000000000000", 31496 => "0000000000000000", 31497 => "0000000000000000", 31498 => "0000000000000000", 31499 => "0000000000000000", 31500 => "0000000000000000", 31501 => "0000000000000000", 31502 => "0000000000000000", 31503 => "0000000000000000", 31504 => "0000000000000000", 31505 => "0000000000000000", 31506 => "0000000000000000", 31507 => "0000000000000000", 31508 => "0000000000000000", 31509 => "0000000000000000", 31510 => "0000000000000000", 31511 => "0000000000000000", 31512 => "0000000000000000", 31513 => "0000000000000000", 31514 => "0000000000000000", 31515 => "0000000000000000", 31516 => "0000000000000000", 31517 => "0000000000000000", 31518 => "0000000000000000", 31519 => "0000000000000000", 31520 => "0000000000000000", 31521 => "0000000000000000", 31522 => "0000000000000000", 31523 => "0000000000000000", 31524 => "0000000000000000", 31525 => "0000000000000000", 31526 => "0000000000000000", 31527 => "0000000000000000", 31528 => "0000000000000000", 31529 => "0000000000000000", 31530 => "0000000000000000", 31531 => "0000000000000000", 31532 => "0000000000000000", 31533 => "0000000000000000", 31534 => "0000000000000000", 31535 => "0000000000000000", 31536 => "0000000000000000", 31537 => "0000000000000000", 31538 => "0000000000000000", 31539 => "0000000000000000", 31540 => "0000000000000000", 31541 => "0000000000000000", 31542 => "0000000000000000", 31543 => "0000000000000000", 31544 => "0000000000000000", 31545 => "0000000000000000", 31546 => "0000000000000000", 31547 => "0000000000000000", 31548 => "0000000000000000", 31549 => "0000000000000000", 31550 => "0000000000000000", 31551 => "0000000000000000", 31552 => "0000000000000000", 31553 => "0000000000000000", 31554 => "0000000000000000", 31555 => "0000000000000000", 31556 => "0000000000000000", 31557 => "0000000000000000", 31558 => "0000000000000000", 31559 => "0000000000000000", 31560 => "0000000000000000", 31561 => "0000000000000000", 31562 => "0000000000000000", 31563 => "0000000000000000", 31564 => "0000000000000000", 31565 => "0000000000000000", 31566 => "0000000000000000", 31567 => "0000000000000000", 31568 => "0000000000000000", 31569 => "0000000000000000", 31570 => "0000000000000000", 31571 => "0000000000000000", 31572 => "0000000000000000", 31573 => "0000000000000000", 31574 => "0000000000000000", 31575 => "0000000000000000", 31576 => "0000000000000000", 31577 => "0000000000000000", 31578 => "0000000000000000", 31579 => "0000000000000000", 31580 => "0000000000000000", 31581 => "0000000000000000", 31582 => "0000000000000000", 31583 => "0000000000000000", 31584 => "0000000000000000", 31585 => "0000000000000000", 31586 => "0000000000000000", 31587 => "0000000000000000", 31588 => "0000000000000000", 31589 => "0000000000000000", 31590 => "0000000000000000", 31591 => "0000000000000000", 31592 => "0000000000000000", 31593 => "0000000000000000", 31594 => "0000000000000000", 31595 => "0000000000000000", 31596 => "0000000000000000", 31597 => "0000000000000000", 31598 => "0000000000000000", 31599 => "0000000000000000", 31600 => "0000000000000000", 31601 => "0000000000000000", 31602 => "0000000000000000", 31603 => "0000000000000000", 31604 => "0000000000000000", 31605 => "0000000000000000", 31606 => "0000000000000000", 31607 => "0000000000000000", 31608 => "0000000000000000", 31609 => "0000000000000000", 31610 => "0000000000000000", 31611 => "0000000000000000", 31612 => "0000000000000000", 31613 => "0000000000000000", 31614 => "0000000000000000", 31615 => "0000000000000000", 31616 => "0000000000000000", 31617 => "0000000000000000", 31618 => "0000000000000000", 31619 => "0000000000000000", 31620 => "0000000000000000", 31621 => "0000000000000000", 31622 => "0000000000000000", 31623 => "0000000000000000", 31624 => "0000000000000000", 31625 => "0000000000000000", 31626 => "0000000000000000", 31627 => "0000000000000000", 31628 => "0000000000000000", 31629 => "0000000000000000", 31630 => "0000000000000000", 31631 => "0000000000000000", 31632 => "0000000000000000", 31633 => "0000000000000000", 31634 => "0000000000000000", 31635 => "0000000000000000", 31636 => "0000000000000000", 31637 => "0000000000000000", 31638 => "0000000000000000", 31639 => "0000000000000000", 31640 => "0000000000000000", 31641 => "0000000000000000", 31642 => "0000000000000000", 31643 => "0000000000000000", 31644 => "0000000000000000", 31645 => "0000000000000000", 31646 => "0000000000000000", 31647 => "0000000000000000", 31648 => "0000000000000000", 31649 => "0000000000000000", 31650 => "0000000000000000", 31651 => "0000000000000000", 31652 => "0000000000000000", 31653 => "0000000000000000", 31654 => "0000000000000000", 31655 => "0000000000000000", 31656 => "0000000000000000", 31657 => "0000000000000000", 31658 => "0000000000000000", 31659 => "0000000000000000", 31660 => "0000000000000000", 31661 => "0000000000000000", 31662 => "0000000000000000", 31663 => "0000000000000000", 31664 => "0000000000000000", 31665 => "0000000000000000", 31666 => "0000000000000000", 31667 => "0000000000000000", 31668 => "0000000000000000", 31669 => "0000000000000000", 31670 => "0000000000000000", 31671 => "0000000000000000", 31672 => "0000000000000000", 31673 => "0000000000000000", 31674 => "0000000000000000", 31675 => "0000000000000000", 31676 => "0000000000000000", 31677 => "0000000000000000", 31678 => "0000000000000000", 31679 => "0000000000000000", 31680 => "0000000000000000", 31681 => "0000000000000000", 31682 => "0000000000000000", 31683 => "0000000000000000", 31684 => "0000000000000000", 31685 => "0000000000000000", 31686 => "0000000000000000", 31687 => "0000000000000000", 31688 => "0000000000000000", 31689 => "0000000000000000", 31690 => "0000000000000000", 31691 => "0000000000000000", 31692 => "0000000000000000", 31693 => "0000000000000000", 31694 => "0000000000000000", 31695 => "0000000000000000", 31696 => "0000000000000000", 31697 => "0000000000000000", 31698 => "0000000000000000", 31699 => "0000000000000000", 31700 => "0000000000000000", 31701 => "0000000000000000", 31702 => "0000000000000000", 31703 => "0000000000000000", 31704 => "0000000000000000", 31705 => "0000000000000000", 31706 => "0000000000000000", 31707 => "0000000000000000", 31708 => "0000000000000000", 31709 => "0000000000000000", 31710 => "0000000000000000", 31711 => "0000000000000000", 31712 => "0000000000000000", 31713 => "0000000000000000", 31714 => "0000000000000000", 31715 => "0000000000000000", 31716 => "0000000000000000", 31717 => "0000000000000000", 31718 => "0000000000000000", 31719 => "0000000000000000", 31720 => "0000000000000000", 31721 => "0000000000000000", 31722 => "0000000000000000", 31723 => "0000000000000000", 31724 => "0000000000000000", 31725 => "0000000000000000", 31726 => "0000000000000000", 31727 => "0000000000000000", 31728 => "0000000000000000", 31729 => "0000000000000000", 31730 => "0000000000000000", 31731 => "0000000000000000", 31732 => "0000000000000000", 31733 => "0000000000000000", 31734 => "0000000000000000", 31735 => "0000000000000000", 31736 => "0000000000000000", 31737 => "0000000000000000", 31738 => "0000000000000000", 31739 => "0000000000000000", 31740 => "0000000000000000", 31741 => "0000000000000000", 31742 => "0000000000000000", 31743 => "0000000000000000", 31744 => "0000000000000000", 31745 => "0000000000000000", 31746 => "0000000000000000", 31747 => "0000000000000000", 31748 => "0000000000000000", 31749 => "0000000000000000", 31750 => "0000000000000000", 31751 => "0000000000000000", 31752 => "0000000000000000", 31753 => "0000000000000000", 31754 => "0000000000000000", 31755 => "0000000000000000", 31756 => "0000000000000000", 31757 => "0000000000000000", 31758 => "0000000000000000", 31759 => "0000000000000000", 31760 => "0000000000000000", 31761 => "0000000000000000", 31762 => "0000000000000000", 31763 => "0000000000000000", 31764 => "0000000000000000", 31765 => "0000000000000000", 31766 => "0000000000000000", 31767 => "0000000000000000", 31768 => "0000000000000000", 31769 => "0000000000000000", 31770 => "0000000000000000", 31771 => "0000000000000000", 31772 => "0000000000000000", 31773 => "0000000000000000", 31774 => "0000000000000000", 31775 => "0000000000000000", 31776 => "0000000000000000", 31777 => "0000000000000000", 31778 => "0000000000000000", 31779 => "0000000000000000", 31780 => "0000000000000000", 31781 => "0000000000000000", 31782 => "0000000000000000", 31783 => "0000000000000000", 31784 => "0000000000000000", 31785 => "0000000000000000", 31786 => "0000000000000000", 31787 => "0000000000000000", 31788 => "0000000000000000", 31789 => "0000000000000000", 31790 => "0000000000000000", 31791 => "0000000000000000", 31792 => "0000000000000000", 31793 => "0000000000000000", 31794 => "0000000000000000", 31795 => "0000000000000000", 31796 => "0000000000000000", 31797 => "0000000000000000", 31798 => "0000000000000000", 31799 => "0000000000000000", 31800 => "0000000000000000", 31801 => "0000000000000000", 31802 => "0000000000000000", 31803 => "0000000000000000", 31804 => "0000000000000000", 31805 => "0000000000000000", 31806 => "0000000000000000", 31807 => "0000000000000000", 31808 => "0000000000000000", 31809 => "0000000000000000", 31810 => "0000000000000000", 31811 => "0000000000000000", 31812 => "0000000000000000", 31813 => "0000000000000000", 31814 => "0000000000000000", 31815 => "0000000000000000", 31816 => "0000000000000000", 31817 => "0000000000000000", 31818 => "0000000000000000", 31819 => "0000000000000000", 31820 => "0000000000000000", 31821 => "0000000000000000", 31822 => "0000000000000000", 31823 => "0000000000000000", 31824 => "0000000000000000", 31825 => "0000000000000000", 31826 => "0000000000000000", 31827 => "0000000000000000", 31828 => "0000000000000000", 31829 => "0000000000000000", 31830 => "0000000000000000", 31831 => "0000000000000000", 31832 => "0000000000000000", 31833 => "0000000000000000", 31834 => "0000000000000000", 31835 => "0000000000000000", 31836 => "0000000000000000", 31837 => "0000000000000000", 31838 => "0000000000000000", 31839 => "0000000000000000", 31840 => "0000000000000000", 31841 => "0000000000000000", 31842 => "0000000000000000", 31843 => "0000000000000000", 31844 => "0000000000000000", 31845 => "0000000000000000", 31846 => "0000000000000000", 31847 => "0000000000000000", 31848 => "0000000000000000", 31849 => "0000000000000000", 31850 => "0000000000000000", 31851 => "0000000000000000", 31852 => "0000000000000000", 31853 => "0000000000000000", 31854 => "0000000000000000", 31855 => "0000000000000000", 31856 => "0000000000000000", 31857 => "0000000000000000", 31858 => "0000000000000000", 31859 => "0000000000000000", 31860 => "0000000000000000", 31861 => "0000000000000000", 31862 => "0000000000000000", 31863 => "0000000000000000", 31864 => "0000000000000000", 31865 => "0000000000000000", 31866 => "0000000000000000", 31867 => "0000000000000000", 31868 => "0000000000000000", 31869 => "0000000000000000", 31870 => "0000000000000000", 31871 => "0000000000000000", 31872 => "0000000000000000", 31873 => "0000000000000000", 31874 => "0000000000000000", 31875 => "0000000000000000", 31876 => "0000000000000000", 31877 => "0000000000000000", 31878 => "0000000000000000", 31879 => "0000000000000000", 31880 => "0000000000000000", 31881 => "0000000000000000", 31882 => "0000000000000000", 31883 => "0000000000000000", 31884 => "0000000000000000", 31885 => "0000000000000000", 31886 => "0000000000000000", 31887 => "0000000000000000", 31888 => "0000000000000000", 31889 => "0000000000000000", 31890 => "0000000000000000", 31891 => "0000000000000000", 31892 => "0000000000000000", 31893 => "0000000000000000", 31894 => "0000000000000000", 31895 => "0000000000000000", 31896 => "0000000000000000", 31897 => "0000000000000000", 31898 => "0000000000000000", 31899 => "0000000000000000", 31900 => "0000000000000000", 31901 => "0000000000000000", 31902 => "0000000000000000", 31903 => "0000000000000000", 31904 => "0000000000000000", 31905 => "0000000000000000", 31906 => "0000000000000000", 31907 => "0000000000000000", 31908 => "0000000000000000", 31909 => "0000000000000000", 31910 => "0000000000000000", 31911 => "0000000000000000", 31912 => "0000000000000000", 31913 => "0000000000000000", 31914 => "0000000000000000", 31915 => "0000000000000000", 31916 => "0000000000000000", 31917 => "0000000000000000", 31918 => "0000000000000000", 31919 => "0000000000000000", 31920 => "0000000000000000", 31921 => "0000000000000000", 31922 => "0000000000000000", 31923 => "0000000000000000", 31924 => "0000000000000000", 31925 => "0000000000000000", 31926 => "0000000000000000", 31927 => "0000000000000000", 31928 => "0000000000000000", 31929 => "0000000000000000", 31930 => "0000000000000000", 31931 => "0000000000000000", 31932 => "0000000000000000", 31933 => "0000000000000000", 31934 => "0000000000000000", 31935 => "0000000000000000", 31936 => "0000000000000000", 31937 => "0000000000000000", 31938 => "0000000000000000", 31939 => "0000000000000000", 31940 => "0000000000000000", 31941 => "0000000000000000", 31942 => "0000000000000000", 31943 => "0000000000000000", 31944 => "0000000000000000", 31945 => "0000000000000000", 31946 => "0000000000000000", 31947 => "0000000000000000", 31948 => "0000000000000000", 31949 => "0000000000000000", 31950 => "0000000000000000", 31951 => "0000000000000000", 31952 => "0000000000000000", 31953 => "0000000000000000", 31954 => "0000000000000000", 31955 => "0000000000000000", 31956 => "0000000000000000", 31957 => "0000000000000000", 31958 => "0000000000000000", 31959 => "0000000000000000", 31960 => "0000000000000000", 31961 => "0000000000000000", 31962 => "0000000000000000", 31963 => "0000000000000000", 31964 => "0000000000000000", 31965 => "0000000000000000", 31966 => "0000000000000000", 31967 => "0000000000000000", 31968 => "0000000000000000", 31969 => "0000000000000000", 31970 => "0000000000000000", 31971 => "0000000000000000", 31972 => "0000000000000000", 31973 => "0000000000000000", 31974 => "0000000000000000", 31975 => "0000000000000000", 31976 => "0000000000000000", 31977 => "0000000000000000", 31978 => "0000000000000000", 31979 => "0000000000000000", 31980 => "0000000000000000", 31981 => "0000000000000000", 31982 => "0000000000000000", 31983 => "0000000000000000", 31984 => "0000000000000000", 31985 => "0000000000000000", 31986 => "0000000000000000", 31987 => "0000000000000000", 31988 => "0000000000000000", 31989 => "0000000000000000", 31990 => "0000000000000000", 31991 => "0000000000000000", 31992 => "0000000000000000", 31993 => "0000000000000000", 31994 => "0000000000000000", 31995 => "0000000000000000", 31996 => "0000000000000000", 31997 => "0000000000000000", 31998 => "0000000000000000", 31999 => "0000000000000000", 32000 => "0000000000000000", 32001 => "0000000000000000", 32002 => "0000000000000000", 32003 => "0000000000000000", 32004 => "0000000000000000", 32005 => "0000000000000000", 32006 => "0000000000000000", 32007 => "0000000000000000", 32008 => "0000000000000000", 32009 => "0000000000000000", 32010 => "0000000000000000", 32011 => "0000000000000000", 32012 => "0000000000000000", 32013 => "0000000000000000", 32014 => "0000000000000000", 32015 => "0000000000000000", 32016 => "0000000000000000", 32017 => "0000000000000000", 32018 => "0000000000000000", 32019 => "0000000000000000", 32020 => "0000000000000000", 32021 => "0000000000000000", 32022 => "0000000000000000", 32023 => "0000000000000000", 32024 => "0000000000000000", 32025 => "0000000000000000", 32026 => "0000000000000000", 32027 => "0000000000000000", 32028 => "0000000000000000", 32029 => "0000000000000000", 32030 => "0000000000000000", 32031 => "0000000000000000", 32032 => "0000000000000000", 32033 => "0000000000000000", 32034 => "0000000000000000", 32035 => "0000000000000000", 32036 => "0000000000000000", 32037 => "0000000000000000", 32038 => "0000000000000000", 32039 => "0000000000000000", 32040 => "0000000000000000", 32041 => "0000000000000000", 32042 => "0000000000000000", 32043 => "0000000000000000", 32044 => "0000000000000000", 32045 => "0000000000000000", 32046 => "0000000000000000", 32047 => "0000000000000000", 32048 => "0000000000000000", 32049 => "0000000000000000", 32050 => "0000000000000000", 32051 => "0000000000000000", 32052 => "0000000000000000", 32053 => "0000000000000000", 32054 => "0000000000000000", 32055 => "0000000000000000", 32056 => "0000000000000000", 32057 => "0000000000000000", 32058 => "0000000000000000", 32059 => "0000000000000000", 32060 => "0000000000000000", 32061 => "0000000000000000", 32062 => "0000000000000000", 32063 => "0000000000000000", 32064 => "0000000000000000", 32065 => "0000000000000000", 32066 => "0000000000000000", 32067 => "0000000000000000", 32068 => "0000000000000000", 32069 => "0000000000000000", 32070 => "0000000000000000", 32071 => "0000000000000000", 32072 => "0000000000000000", 32073 => "0000000000000000", 32074 => "0000000000000000", 32075 => "0000000000000000", 32076 => "0000000000000000", 32077 => "0000000000000000", 32078 => "0000000000000000", 32079 => "0000000000000000", 32080 => "0000000000000000", 32081 => "0000000000000000", 32082 => "0000000000000000", 32083 => "0000000000000000", 32084 => "0000000000000000", 32085 => "0000000000000000", 32086 => "0000000000000000", 32087 => "0000000000000000", 32088 => "0000000000000000", 32089 => "0000000000000000", 32090 => "0000000000000000", 32091 => "0000000000000000", 32092 => "0000000000000000", 32093 => "0000000000000000", 32094 => "0000000000000000", 32095 => "0000000000000000", 32096 => "0000000000000000", 32097 => "0000000000000000", 32098 => "0000000000000000", 32099 => "0000000000000000", 32100 => "0000000000000000", 32101 => "0000000000000000", 32102 => "0000000000000000", 32103 => "0000000000000000", 32104 => "0000000000000000", 32105 => "0000000000000000", 32106 => "0000000000000000", 32107 => "0000000000000000", 32108 => "0000000000000000", 32109 => "0000000000000000", 32110 => "0000000000000000", 32111 => "0000000000000000", 32112 => "0000000000000000", 32113 => "0000000000000000", 32114 => "0000000000000000", 32115 => "0000000000000000", 32116 => "0000000000000000", 32117 => "0000000000000000", 32118 => "0000000000000000", 32119 => "0000000000000000", 32120 => "0000000000000000", 32121 => "0000000000000000", 32122 => "0000000000000000", 32123 => "0000000000000000", 32124 => "0000000000000000", 32125 => "0000000000000000", 32126 => "0000000000000000", 32127 => "0000000000000000", 32128 => "0000000000000000", 32129 => "0000000000000000", 32130 => "0000000000000000", 32131 => "0000000000000000", 32132 => "0000000000000000", 32133 => "0000000000000000", 32134 => "0000000000000000", 32135 => "0000000000000000", 32136 => "0000000000000000", 32137 => "0000000000000000", 32138 => "0000000000000000", 32139 => "0000000000000000", 32140 => "0000000000000000", 32141 => "0000000000000000", 32142 => "0000000000000000", 32143 => "0000000000000000", 32144 => "0000000000000000", 32145 => "0000000000000000", 32146 => "0000000000000000", 32147 => "0000000000000000", 32148 => "0000000000000000", 32149 => "0000000000000000", 32150 => "0000000000000000", 32151 => "0000000000000000", 32152 => "0000000000000000", 32153 => "0000000000000000", 32154 => "0000000000000000", 32155 => "0000000000000000", 32156 => "0000000000000000", 32157 => "0000000000000000", 32158 => "0000000000000000", 32159 => "0000000000000000", 32160 => "0000000000000000", 32161 => "0000000000000000", 32162 => "0000000000000000", 32163 => "0000000000000000", 32164 => "0000000000000000", 32165 => "0000000000000000", 32166 => "0000000000000000", 32167 => "0000000000000000", 32168 => "0000000000000000", 32169 => "0000000000000000", 32170 => "0000000000000000", 32171 => "0000000000000000", 32172 => "0000000000000000", 32173 => "0000000000000000", 32174 => "0000000000000000", 32175 => "0000000000000000", 32176 => "0000000000000000", 32177 => "0000000000000000", 32178 => "0000000000000000", 32179 => "0000000000000000", 32180 => "0000000000000000", 32181 => "0000000000000000", 32182 => "0000000000000000", 32183 => "0000000000000000", 32184 => "0000000000000000", 32185 => "0000000000000000", 32186 => "0000000000000000", 32187 => "0000000000000000", 32188 => "0000000000000000", 32189 => "0000000000000000", 32190 => "0000000000000000", 32191 => "0000000000000000", 32192 => "0000000000000000", 32193 => "0000000000000000", 32194 => "0000000000000000", 32195 => "0000000000000000", 32196 => "0000000000000000", 32197 => "0000000000000000", 32198 => "0000000000000000", 32199 => "0000000000000000", 32200 => "0000000000000000", 32201 => "0000000000000000", 32202 => "0000000000000000", 32203 => "0000000000000000", 32204 => "0000000000000000", 32205 => "0000000000000000", 32206 => "0000000000000000", 32207 => "0000000000000000", 32208 => "0000000000000000", 32209 => "0000000000000000", 32210 => "0000000000000000", 32211 => "0000000000000000", 32212 => "0000000000000000", 32213 => "0000000000000000", 32214 => "0000000000000000", 32215 => "0000000000000000", 32216 => "0000000000000000", 32217 => "0000000000000000", 32218 => "0000000000000000", 32219 => "0000000000000000", 32220 => "0000000000000000", 32221 => "0000000000000000", 32222 => "0000000000000000", 32223 => "0000000000000000", 32224 => "0000000000000000", 32225 => "0000000000000000", 32226 => "0000000000000000", 32227 => "0000000000000000", 32228 => "0000000000000000", 32229 => "0000000000000000", 32230 => "0000000000000000", 32231 => "0000000000000000", 32232 => "0000000000000000", 32233 => "0000000000000000", 32234 => "0000000000000000", 32235 => "0000000000000000", 32236 => "0000000000000000", 32237 => "0000000000000000", 32238 => "0000000000000000", 32239 => "0000000000000000", 32240 => "0000000000000000", 32241 => "0000000000000000", 32242 => "0000000000000000", 32243 => "0000000000000000", 32244 => "0000000000000000", 32245 => "0000000000000000", 32246 => "0000000000000000", 32247 => "0000000000000000", 32248 => "0000000000000000", 32249 => "0000000000000000", 32250 => "0000000000000000", 32251 => "0000000000000000", 32252 => "0000000000000000", 32253 => "0000000000000000", 32254 => "0000000000000000", 32255 => "0000000000000000", 32256 => "0000000000000000", 32257 => "0000000000000000", 32258 => "0000000000000000", 32259 => "0000000000000000", 32260 => "0000000000000000", 32261 => "0000000000000000", 32262 => "0000000000000000", 32263 => "0000000000000000", 32264 => "0000000000000000", 32265 => "0000000000000000", 32266 => "0000000000000000", 32267 => "0000000000000000", 32268 => "0000000000000000", 32269 => "0000000000000000", 32270 => "0000000000000000", 32271 => "0000000000000000", 32272 => "0000000000000000", 32273 => "0000000000000000", 32274 => "0000000000000000", 32275 => "0000000000000000", 32276 => "0000000000000000", 32277 => "0000000000000000", 32278 => "0000000000000000", 32279 => "0000000000000000", 32280 => "0000000000000000", 32281 => "0000000000000000", 32282 => "0000000000000000", 32283 => "0000000000000000", 32284 => "0000000000000000", 32285 => "0000000000000000", 32286 => "0000000000000000", 32287 => "0000000000000000", 32288 => "0000000000000000", 32289 => "0000000000000000", 32290 => "0000000000000000", 32291 => "0000000000000000", 32292 => "0000000000000000", 32293 => "0000000000000000", 32294 => "0000000000000000", 32295 => "0000000000000000", 32296 => "0000000000000000", 32297 => "0000000000000000", 32298 => "0000000000000000", 32299 => "0000000000000000", 32300 => "0000000000000000", 32301 => "0000000000000000", 32302 => "0000000000000000", 32303 => "0000000000000000", 32304 => "0000000000000000", 32305 => "0000000000000000", 32306 => "0000000000000000", 32307 => "0000000000000000", 32308 => "0000000000000000", 32309 => "0000000000000000", 32310 => "0000000000000000", 32311 => "0000000000000000", 32312 => "0000000000000000", 32313 => "0000000000000000", 32314 => "0000000000000000", 32315 => "0000000000000000", 32316 => "0000000000000000", 32317 => "0000000000000000", 32318 => "0000000000000000", 32319 => "0000000000000000", 32320 => "0000000000000000", 32321 => "0000000000000000", 32322 => "0000000000000000", 32323 => "0000000000000000", 32324 => "0000000000000000", 32325 => "0000000000000000", 32326 => "0000000000000000", 32327 => "0000000000000000", 32328 => "0000000000000000", 32329 => "0000000000000000", 32330 => "0000000000000000", 32331 => "0000000000000000", 32332 => "0000000000000000", 32333 => "0000000000000000", 32334 => "0000000000000000", 32335 => "0000000000000000", 32336 => "0000000000000000", 32337 => "0000000000000000", 32338 => "0000000000000000", 32339 => "0000000000000000", 32340 => "0000000000000000", 32341 => "0000000000000000", 32342 => "0000000000000000", 32343 => "0000000000000000", 32344 => "0000000000000000", 32345 => "0000000000000000", 32346 => "0000000000000000", 32347 => "0000000000000000", 32348 => "0000000000000000", 32349 => "0000000000000000", 32350 => "0000000000000000", 32351 => "0000000000000000", 32352 => "0000000000000000", 32353 => "0000000000000000", 32354 => "0000000000000000", 32355 => "0000000000000000", 32356 => "0000000000000000", 32357 => "0000000000000000", 32358 => "0000000000000000", 32359 => "0000000000000000", 32360 => "0000000000000000", 32361 => "0000000000000000", 32362 => "0000000000000000", 32363 => "0000000000000000", 32364 => "0000000000000000", 32365 => "0000000000000000", 32366 => "0000000000000000", 32367 => "0000000000000000", 32368 => "0000000000000000", 32369 => "0000000000000000", 32370 => "0000000000000000", 32371 => "0000000000000000", 32372 => "0000000000000000", 32373 => "0000000000000000", 32374 => "0000000000000000", 32375 => "0000000000000000", 32376 => "0000000000000000", 32377 => "0000000000000000", 32378 => "0000000000000000", 32379 => "0000000000000000", 32380 => "0000000000000000", 32381 => "0000000000000000", 32382 => "0000000000000000", 32383 => "0000000000000000", 32384 => "0000000000000000", 32385 => "0000000000000000", 32386 => "0000000000000000", 32387 => "0000000000000000", 32388 => "0000000000000000", 32389 => "0000000000000000", 32390 => "0000000000000000", 32391 => "0000000000000000", 32392 => "0000000000000000", 32393 => "0000000000000000", 32394 => "0000000000000000", 32395 => "0000000000000000", 32396 => "0000000000000000", 32397 => "0000000000000000", 32398 => "0000000000000000", 32399 => "0000000000000000", 32400 => "0000000000000000", 32401 => "0000000000000000", 32402 => "0000000000000000", 32403 => "0000000000000000", 32404 => "0000000000000000", 32405 => "0000000000000000", 32406 => "0000000000000000", 32407 => "0000000000000000", 32408 => "0000000000000000", 32409 => "0000000000000000", 32410 => "0000000000000000", 32411 => "0000000000000000", 32412 => "0000000000000000", 32413 => "0000000000000000", 32414 => "0000000000000000", 32415 => "0000000000000000", 32416 => "0000000000000000", 32417 => "0000000000000000", 32418 => "0000000000000000", 32419 => "0000000000000000", 32420 => "0000000000000000", 32421 => "0000000000000000", 32422 => "0000000000000000", 32423 => "0000000000000000", 32424 => "0000000000000000", 32425 => "0000000000000000", 32426 => "0000000000000000", 32427 => "0000000000000000", 32428 => "0000000000000000", 32429 => "0000000000000000", 32430 => "0000000000000000", 32431 => "0000000000000000", 32432 => "0000000000000000", 32433 => "0000000000000000", 32434 => "0000000000000000", 32435 => "0000000000000000", 32436 => "0000000000000000", 32437 => "0000000000000000", 32438 => "0000000000000000", 32439 => "0000000000000000", 32440 => "0000000000000000", 32441 => "0000000000000000", 32442 => "0000000000000000", 32443 => "0000000000000000", 32444 => "0000000000000000", 32445 => "0000000000000000", 32446 => "0000000000000000", 32447 => "0000000000000000", 32448 => "0000000000000000", 32449 => "0000000000000000", 32450 => "0000000000000000", 32451 => "0000000000000000", 32452 => "0000000000000000", 32453 => "0000000000000000", 32454 => "0000000000000000", 32455 => "0000000000000000", 32456 => "0000000000000000", 32457 => "0000000000000000", 32458 => "0000000000000000", 32459 => "0000000000000000", 32460 => "0000000000000000", 32461 => "0000000000000000", 32462 => "0000000000000000", 32463 => "0000000000000000", 32464 => "0000000000000000", 32465 => "0000000000000000", 32466 => "0000000000000000", 32467 => "0000000000000000", 32468 => "0000000000000000", 32469 => "0000000000000000", 32470 => "0000000000000000", 32471 => "0000000000000000", 32472 => "0000000000000000", 32473 => "0000000000000000", 32474 => "0000000000000000", 32475 => "0000000000000000", 32476 => "0000000000000000", 32477 => "0000000000000000", 32478 => "0000000000000000", 32479 => "0000000000000000", 32480 => "0000000000000000", 32481 => "0000000000000000", 32482 => "0000000000000000", 32483 => "0000000000000000", 32484 => "0000000000000000", 32485 => "0000000000000000", 32486 => "0000000000000000", 32487 => "0000000000000000", 32488 => "0000000000000000", 32489 => "0000000000000000", 32490 => "0000000000000000", 32491 => "0000000000000000", 32492 => "0000000000000000", 32493 => "0000000000000000", 32494 => "0000000000000000", 32495 => "0000000000000000", 32496 => "0000000000000000", 32497 => "0000000000000000", 32498 => "0000000000000000", 32499 => "0000000000000000", 32500 => "0000000000000000", 32501 => "0000000000000000", 32502 => "0000000000000000", 32503 => "0000000000000000", 32504 => "0000000000000000", 32505 => "0000000000000000", 32506 => "0000000000000000", 32507 => "0000000000000000", 32508 => "0000000000000000", 32509 => "0000000000000000", 32510 => "0000000000000000", 32511 => "0000000000000000", 32512 => "0000000000000000", 32513 => "0000000000000000", 32514 => "0000000000000000", 32515 => "0000000000000000", 32516 => "0000000000000000", 32517 => "0000000000000000", 32518 => "0000000000000000", 32519 => "0000000000000000", 32520 => "0000000000000000", 32521 => "0000000000000000", 32522 => "0000000000000000", 32523 => "0000000000000000", 32524 => "0000000000000000", 32525 => "0000000000000000", 32526 => "0000000000000000", 32527 => "0000000000000000", 32528 => "0000000000000000", 32529 => "0000000000000000", 32530 => "0000000000000000", 32531 => "0000000000000000", 32532 => "0000000000000000", 32533 => "0000000000000000", 32534 => "0000000000000000", 32535 => "0000000000000000", 32536 => "0000000000000000", 32537 => "0000000000000000", 32538 => "0000000000000000", 32539 => "0000000000000000", 32540 => "0000000000000000", 32541 => "0000000000000000", 32542 => "0000000000000000", 32543 => "0000000000000000", 32544 => "0000000000000000", 32545 => "0000000000000000", 32546 => "0000000000000000", 32547 => "0000000000000000", 32548 => "0000000000000000", 32549 => "0000000000000000", 32550 => "0000000000000000", 32551 => "0000000000000000", 32552 => "0000000000000000", 32553 => "0000000000000000", 32554 => "0000000000000000", 32555 => "0000000000000000", 32556 => "0000000000000000", 32557 => "0000000000000000", 32558 => "0000000000000000", 32559 => "0000000000000000", 32560 => "0000000000000000", 32561 => "0000000000000000", 32562 => "0000000000000000", 32563 => "0000000000000000", 32564 => "0000000000000000", 32565 => "0000000000000000", 32566 => "0000000000000000", 32567 => "0000000000000000", 32568 => "0000000000000000", 32569 => "0000000000000000", 32570 => "0000000000000000", 32571 => "0000000000000000", 32572 => "0000000000000000", 32573 => "0000000000000000", 32574 => "0000000000000000", 32575 => "0000000000000000", 32576 => "0000000000000000", 32577 => "0000000000000000", 32578 => "0000000000000000", 32579 => "0000000000000000", 32580 => "0000000000000000", 32581 => "0000000000000000", 32582 => "0000000000000000", 32583 => "0000000000000000", 32584 => "0000000000000000", 32585 => "0000000000000000", 32586 => "0000000000000000", 32587 => "0000000000000000", 32588 => "0000000000000000", 32589 => "0000000000000000", 32590 => "0000000000000000", 32591 => "0000000000000000", 32592 => "0000000000000000", 32593 => "0000000000000000", 32594 => "0000000000000000", 32595 => "0000000000000000", 32596 => "0000000000000000", 32597 => "0000000000000000", 32598 => "0000000000000000", 32599 => "0000000000000000", 32600 => "0000000000000000", 32601 => "0000000000000000", 32602 => "0000000000000000", 32603 => "0000000000000000", 32604 => "0000000000000000", 32605 => "0000000000000000", 32606 => "0000000000000000", 32607 => "0000000000000000", 32608 => "0000000000000000", 32609 => "0000000000000000", 32610 => "0000000000000000", 32611 => "0000000000000000", 32612 => "0000000000000000", 32613 => "0000000000000000", 32614 => "0000000000000000", 32615 => "0000000000000000", 32616 => "0000000000000000", 32617 => "0000000000000000", 32618 => "0000000000000000", 32619 => "0000000000000000", 32620 => "0000000000000000", 32621 => "0000000000000000", 32622 => "0000000000000000", 32623 => "0000000000000000", 32624 => "0000000000000000", 32625 => "0000000000000000", 32626 => "0000000000000000", 32627 => "0000000000000000", 32628 => "0000000000000000", 32629 => "0000000000000000", 32630 => "0000000000000000", 32631 => "0000000000000000", 32632 => "0000000000000000", 32633 => "0000000000000000", 32634 => "0000000000000000", 32635 => "0000000000000000", 32636 => "0000000000000000", 32637 => "0000000000000000", 32638 => "0000000000000000", 32639 => "0000000000000000", 32640 => "0000000000000000", 32641 => "0000000000000000", 32642 => "0000000000000000", 32643 => "0000000000000000", 32644 => "0000000000000000", 32645 => "0000000000000000", 32646 => "0000000000000000", 32647 => "0000000000000000", 32648 => "0000000000000000", 32649 => "0000000000000000", 32650 => "0000000000000000", 32651 => "0000000000000000", 32652 => "0000000000000000", 32653 => "0000000000000000", 32654 => "0000000000000000", 32655 => "0000000000000000", 32656 => "0000000000000000", 32657 => "0000000000000000", 32658 => "0000000000000000", 32659 => "0000000000000000", 32660 => "0000000000000000", 32661 => "0000000000000000", 32662 => "0000000000000000", 32663 => "0000000000000000", 32664 => "0000000000000000", 32665 => "0000000000000000", 32666 => "0000000000000000", 32667 => "0000000000000000", 32668 => "0000000000000000", 32669 => "0000000000000000", 32670 => "0000000000000000", 32671 => "0000000000000000", 32672 => "0000000000000000", 32673 => "0000000000000000", 32674 => "0000000000000000", 32675 => "0000000000000000", 32676 => "0000000000000000", 32677 => "0000000000000000", 32678 => "0000000000000000", 32679 => "0000000000000000", 32680 => "0000000000000000", 32681 => "0000000000000000", 32682 => "0000000000000000", 32683 => "0000000000000000", 32684 => "0000000000000000", 32685 => "0000000000000000", 32686 => "0000000000000000", 32687 => "0000000000000000", 32688 => "0000000000000000", 32689 => "0000000000000000", 32690 => "0000000000000000", 32691 => "0000000000000000", 32692 => "0000000000000000", 32693 => "0000000000000000", 32694 => "0000000000000000", 32695 => "0000000000000000", 32696 => "0000000000000000", 32697 => "0000000000000000", 32698 => "0000000000000000", 32699 => "0000000000000000", 32700 => "0000000000000000", 32701 => "0000000000000000", 32702 => "0000000000000000", 32703 => "0000000000000000", 32704 => "0000000000000000", 32705 => "0000000000000000", 32706 => "0000000000000000", 32707 => "0000000000000000", 32708 => "0000000000000000", 32709 => "0000000000000000", 32710 => "0000000000000000", 32711 => "0000000000000000", 32712 => "0000000000000000", 32713 => "0000000000000000", 32714 => "0000000000000000", 32715 => "0000000000000000", 32716 => "0000000000000000", 32717 => "0000000000000000", 32718 => "0000000000000000", 32719 => "0000000000000000", 32720 => "0000000000000000", 32721 => "0000000000000000", 32722 => "0000000000000000", 32723 => "0000000000000000", 32724 => "0000000000000000", 32725 => "0000000000000000", 32726 => "0000000000000000", 32727 => "0000000000000000", 32728 => "0000000000000000", 32729 => "0000000000000000", 32730 => "0000000000000000", 32731 => "0000000000000000", 32732 => "0000000000000000", 32733 => "0000000000000000", 32734 => "0000000000000000", 32735 => "0000000000000000", 32736 => "0000000000000000", 32737 => "0000000000000000", 32738 => "0000000000000000", 32739 => "0000000000000000", 32740 => "0000000000000000", 32741 => "0000000000000000", 32742 => "0000000000000000", 32743 => "0000000000000000", 32744 => "0000000000000000", 32745 => "0000000000000000", 32746 => "0000000000000000", 32747 => "0000000000000000", 32748 => "0000000000000000", 32749 => "0000000000000000", 32750 => "0000000000000000", 32751 => "0000000000000000", 32752 => "0000000000000000", 32753 => "0000000000000000", 32754 => "0000000000000000", 32755 => "0000000000000000", 32756 => "0000000000000000", 32757 => "0000000000000000", 32758 => "0000000000000000", 32759 => "0000000000000000", 32760 => "0000000000000000", 32761 => "0000000000000000", 32762 => "0000000000000000", 32763 => "0000000000000000", 32764 => "0000000000000000", 32765 => "0000000000000000", 32766 => "0000000000000000", 32767 => "0000000000000000");
BEGIN
  data_out <= ROM(to_integer(unsigned(address)));
END ARCHITECTURE;
